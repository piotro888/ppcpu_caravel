* NGSPICE file created from interconnect_inner.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

.subckt interconnect_inner c0_clk c0_dbg_pc[0] c0_dbg_pc[10] c0_dbg_pc[11] c0_dbg_pc[12]
+ c0_dbg_pc[13] c0_dbg_pc[14] c0_dbg_pc[15] c0_dbg_pc[1] c0_dbg_pc[2] c0_dbg_pc[3]
+ c0_dbg_pc[4] c0_dbg_pc[5] c0_dbg_pc[6] c0_dbg_pc[7] c0_dbg_pc[8] c0_dbg_pc[9] c0_dbg_r0[0]
+ c0_dbg_r0[10] c0_dbg_r0[11] c0_dbg_r0[12] c0_dbg_r0[13] c0_dbg_r0[14] c0_dbg_r0[15]
+ c0_dbg_r0[1] c0_dbg_r0[2] c0_dbg_r0[3] c0_dbg_r0[4] c0_dbg_r0[5] c0_dbg_r0[6] c0_dbg_r0[7]
+ c0_dbg_r0[8] c0_dbg_r0[9] c0_disable c0_i_core_int_sreg[0] c0_i_core_int_sreg[10]
+ c0_i_core_int_sreg[11] c0_i_core_int_sreg[12] c0_i_core_int_sreg[13] c0_i_core_int_sreg[14]
+ c0_i_core_int_sreg[15] c0_i_core_int_sreg[1] c0_i_core_int_sreg[2] c0_i_core_int_sreg[3]
+ c0_i_core_int_sreg[4] c0_i_core_int_sreg[5] c0_i_core_int_sreg[6] c0_i_core_int_sreg[7]
+ c0_i_core_int_sreg[8] c0_i_core_int_sreg[9] c0_i_irq c0_i_mc_core_int c0_i_mem_ack
+ c0_i_mem_data[0] c0_i_mem_data[10] c0_i_mem_data[11] c0_i_mem_data[12] c0_i_mem_data[13]
+ c0_i_mem_data[14] c0_i_mem_data[15] c0_i_mem_data[1] c0_i_mem_data[2] c0_i_mem_data[3]
+ c0_i_mem_data[4] c0_i_mem_data[5] c0_i_mem_data[6] c0_i_mem_data[7] c0_i_mem_data[8]
+ c0_i_mem_data[9] c0_i_mem_exception c0_i_req_data[0] c0_i_req_data[10] c0_i_req_data[11]
+ c0_i_req_data[12] c0_i_req_data[13] c0_i_req_data[14] c0_i_req_data[15] c0_i_req_data[16]
+ c0_i_req_data[17] c0_i_req_data[18] c0_i_req_data[19] c0_i_req_data[1] c0_i_req_data[20]
+ c0_i_req_data[21] c0_i_req_data[22] c0_i_req_data[23] c0_i_req_data[24] c0_i_req_data[25]
+ c0_i_req_data[26] c0_i_req_data[27] c0_i_req_data[28] c0_i_req_data[29] c0_i_req_data[2]
+ c0_i_req_data[30] c0_i_req_data[31] c0_i_req_data[3] c0_i_req_data[4] c0_i_req_data[5]
+ c0_i_req_data[6] c0_i_req_data[7] c0_i_req_data[8] c0_i_req_data[9] c0_i_req_data_valid
+ c0_o_c_data_page c0_o_c_instr_long c0_o_c_instr_page c0_o_icache_flush c0_o_instr_long_addr[0]
+ c0_o_instr_long_addr[1] c0_o_instr_long_addr[2] c0_o_instr_long_addr[3] c0_o_instr_long_addr[4]
+ c0_o_instr_long_addr[5] c0_o_instr_long_addr[6] c0_o_instr_long_addr[7] c0_o_mem_addr[0]
+ c0_o_mem_addr[10] c0_o_mem_addr[11] c0_o_mem_addr[12] c0_o_mem_addr[13] c0_o_mem_addr[14]
+ c0_o_mem_addr[15] c0_o_mem_addr[1] c0_o_mem_addr[2] c0_o_mem_addr[3] c0_o_mem_addr[4]
+ c0_o_mem_addr[5] c0_o_mem_addr[6] c0_o_mem_addr[7] c0_o_mem_addr[8] c0_o_mem_addr[9]
+ c0_o_mem_data[0] c0_o_mem_data[10] c0_o_mem_data[11] c0_o_mem_data[12] c0_o_mem_data[13]
+ c0_o_mem_data[14] c0_o_mem_data[15] c0_o_mem_data[1] c0_o_mem_data[2] c0_o_mem_data[3]
+ c0_o_mem_data[4] c0_o_mem_data[5] c0_o_mem_data[6] c0_o_mem_data[7] c0_o_mem_data[8]
+ c0_o_mem_data[9] c0_o_mem_high_addr[0] c0_o_mem_high_addr[1] c0_o_mem_high_addr[2]
+ c0_o_mem_high_addr[3] c0_o_mem_high_addr[4] c0_o_mem_high_addr[5] c0_o_mem_high_addr[6]
+ c0_o_mem_high_addr[7] c0_o_mem_long_mode c0_o_mem_req c0_o_mem_sel[0] c0_o_mem_sel[1]
+ c0_o_mem_we c0_o_req_active c0_o_req_addr[0] c0_o_req_addr[10] c0_o_req_addr[11]
+ c0_o_req_addr[12] c0_o_req_addr[13] c0_o_req_addr[14] c0_o_req_addr[15] c0_o_req_addr[1]
+ c0_o_req_addr[2] c0_o_req_addr[3] c0_o_req_addr[4] c0_o_req_addr[5] c0_o_req_addr[6]
+ c0_o_req_addr[7] c0_o_req_addr[8] c0_o_req_addr[9] c0_o_req_ppl_submit c0_rst c0_sr_bus_addr[0]
+ c0_sr_bus_addr[10] c0_sr_bus_addr[11] c0_sr_bus_addr[12] c0_sr_bus_addr[13] c0_sr_bus_addr[14]
+ c0_sr_bus_addr[15] c0_sr_bus_addr[1] c0_sr_bus_addr[2] c0_sr_bus_addr[3] c0_sr_bus_addr[4]
+ c0_sr_bus_addr[5] c0_sr_bus_addr[6] c0_sr_bus_addr[7] c0_sr_bus_addr[8] c0_sr_bus_addr[9]
+ c0_sr_bus_data_o[0] c0_sr_bus_data_o[10] c0_sr_bus_data_o[11] c0_sr_bus_data_o[12]
+ c0_sr_bus_data_o[13] c0_sr_bus_data_o[14] c0_sr_bus_data_o[15] c0_sr_bus_data_o[1]
+ c0_sr_bus_data_o[2] c0_sr_bus_data_o[3] c0_sr_bus_data_o[4] c0_sr_bus_data_o[5]
+ c0_sr_bus_data_o[6] c0_sr_bus_data_o[7] c0_sr_bus_data_o[8] c0_sr_bus_data_o[9]
+ c0_sr_bus_we c1_clk c1_dbg_pc[0] c1_dbg_pc[10] c1_dbg_pc[11] c1_dbg_pc[12] c1_dbg_pc[13]
+ c1_dbg_pc[14] c1_dbg_pc[15] c1_dbg_pc[1] c1_dbg_pc[2] c1_dbg_pc[3] c1_dbg_pc[4]
+ c1_dbg_pc[5] c1_dbg_pc[6] c1_dbg_pc[7] c1_dbg_pc[8] c1_dbg_pc[9] c1_dbg_r0[0] c1_dbg_r0[10]
+ c1_dbg_r0[11] c1_dbg_r0[12] c1_dbg_r0[13] c1_dbg_r0[14] c1_dbg_r0[15] c1_dbg_r0[1]
+ c1_dbg_r0[2] c1_dbg_r0[3] c1_dbg_r0[4] c1_dbg_r0[5] c1_dbg_r0[6] c1_dbg_r0[7] c1_dbg_r0[8]
+ c1_dbg_r0[9] c1_disable c1_i_core_int_sreg[0] c1_i_core_int_sreg[10] c1_i_core_int_sreg[11]
+ c1_i_core_int_sreg[12] c1_i_core_int_sreg[13] c1_i_core_int_sreg[14] c1_i_core_int_sreg[15]
+ c1_i_core_int_sreg[1] c1_i_core_int_sreg[2] c1_i_core_int_sreg[3] c1_i_core_int_sreg[4]
+ c1_i_core_int_sreg[5] c1_i_core_int_sreg[6] c1_i_core_int_sreg[7] c1_i_core_int_sreg[8]
+ c1_i_core_int_sreg[9] c1_i_irq c1_i_mc_core_int c1_i_mem_ack c1_i_mem_data[0] c1_i_mem_data[10]
+ c1_i_mem_data[11] c1_i_mem_data[12] c1_i_mem_data[13] c1_i_mem_data[14] c1_i_mem_data[15]
+ c1_i_mem_data[1] c1_i_mem_data[2] c1_i_mem_data[3] c1_i_mem_data[4] c1_i_mem_data[5]
+ c1_i_mem_data[6] c1_i_mem_data[7] c1_i_mem_data[8] c1_i_mem_data[9] c1_i_mem_exception
+ c1_i_req_data[0] c1_i_req_data[10] c1_i_req_data[11] c1_i_req_data[12] c1_i_req_data[13]
+ c1_i_req_data[14] c1_i_req_data[15] c1_i_req_data[16] c1_i_req_data[17] c1_i_req_data[18]
+ c1_i_req_data[19] c1_i_req_data[1] c1_i_req_data[20] c1_i_req_data[21] c1_i_req_data[22]
+ c1_i_req_data[23] c1_i_req_data[24] c1_i_req_data[25] c1_i_req_data[26] c1_i_req_data[27]
+ c1_i_req_data[28] c1_i_req_data[29] c1_i_req_data[2] c1_i_req_data[30] c1_i_req_data[31]
+ c1_i_req_data[3] c1_i_req_data[4] c1_i_req_data[5] c1_i_req_data[6] c1_i_req_data[7]
+ c1_i_req_data[8] c1_i_req_data[9] c1_i_req_data_valid c1_o_c_data_page c1_o_c_instr_long
+ c1_o_c_instr_page c1_o_icache_flush c1_o_instr_long_addr[0] c1_o_instr_long_addr[1]
+ c1_o_instr_long_addr[2] c1_o_instr_long_addr[3] c1_o_instr_long_addr[4] c1_o_instr_long_addr[5]
+ c1_o_instr_long_addr[6] c1_o_instr_long_addr[7] c1_o_mem_addr[0] c1_o_mem_addr[10]
+ c1_o_mem_addr[11] c1_o_mem_addr[12] c1_o_mem_addr[13] c1_o_mem_addr[14] c1_o_mem_addr[15]
+ c1_o_mem_addr[1] c1_o_mem_addr[2] c1_o_mem_addr[3] c1_o_mem_addr[4] c1_o_mem_addr[5]
+ c1_o_mem_addr[6] c1_o_mem_addr[7] c1_o_mem_addr[8] c1_o_mem_addr[9] c1_o_mem_data[0]
+ c1_o_mem_data[10] c1_o_mem_data[11] c1_o_mem_data[12] c1_o_mem_data[13] c1_o_mem_data[14]
+ c1_o_mem_data[15] c1_o_mem_data[1] c1_o_mem_data[2] c1_o_mem_data[3] c1_o_mem_data[4]
+ c1_o_mem_data[5] c1_o_mem_data[6] c1_o_mem_data[7] c1_o_mem_data[8] c1_o_mem_data[9]
+ c1_o_mem_high_addr[0] c1_o_mem_high_addr[1] c1_o_mem_high_addr[2] c1_o_mem_high_addr[3]
+ c1_o_mem_high_addr[4] c1_o_mem_high_addr[5] c1_o_mem_high_addr[6] c1_o_mem_high_addr[7]
+ c1_o_mem_long_mode c1_o_mem_req c1_o_mem_sel[0] c1_o_mem_sel[1] c1_o_mem_we c1_o_req_active
+ c1_o_req_addr[0] c1_o_req_addr[10] c1_o_req_addr[11] c1_o_req_addr[12] c1_o_req_addr[13]
+ c1_o_req_addr[14] c1_o_req_addr[15] c1_o_req_addr[1] c1_o_req_addr[2] c1_o_req_addr[3]
+ c1_o_req_addr[4] c1_o_req_addr[5] c1_o_req_addr[6] c1_o_req_addr[7] c1_o_req_addr[8]
+ c1_o_req_addr[9] c1_o_req_ppl_submit c1_rst c1_sr_bus_addr[0] c1_sr_bus_addr[10]
+ c1_sr_bus_addr[11] c1_sr_bus_addr[12] c1_sr_bus_addr[13] c1_sr_bus_addr[14] c1_sr_bus_addr[15]
+ c1_sr_bus_addr[1] c1_sr_bus_addr[2] c1_sr_bus_addr[3] c1_sr_bus_addr[4] c1_sr_bus_addr[5]
+ c1_sr_bus_addr[6] c1_sr_bus_addr[7] c1_sr_bus_addr[8] c1_sr_bus_addr[9] c1_sr_bus_data_o[0]
+ c1_sr_bus_data_o[10] c1_sr_bus_data_o[11] c1_sr_bus_data_o[12] c1_sr_bus_data_o[13]
+ c1_sr_bus_data_o[14] c1_sr_bus_data_o[15] c1_sr_bus_data_o[1] c1_sr_bus_data_o[2]
+ c1_sr_bus_data_o[3] c1_sr_bus_data_o[4] c1_sr_bus_data_o[5] c1_sr_bus_data_o[6]
+ c1_sr_bus_data_o[7] c1_sr_bus_data_o[8] c1_sr_bus_data_o[9] c1_sr_bus_we core_clock
+ core_reset dcache_clk dcache_mem_ack dcache_mem_addr[0] dcache_mem_addr[10] dcache_mem_addr[11]
+ dcache_mem_addr[12] dcache_mem_addr[13] dcache_mem_addr[14] dcache_mem_addr[15]
+ dcache_mem_addr[16] dcache_mem_addr[17] dcache_mem_addr[18] dcache_mem_addr[19]
+ dcache_mem_addr[1] dcache_mem_addr[20] dcache_mem_addr[21] dcache_mem_addr[22] dcache_mem_addr[23]
+ dcache_mem_addr[2] dcache_mem_addr[3] dcache_mem_addr[4] dcache_mem_addr[5] dcache_mem_addr[6]
+ dcache_mem_addr[7] dcache_mem_addr[8] dcache_mem_addr[9] dcache_mem_cache_enable
+ dcache_mem_exception dcache_mem_i_data[0] dcache_mem_i_data[10] dcache_mem_i_data[11]
+ dcache_mem_i_data[12] dcache_mem_i_data[13] dcache_mem_i_data[14] dcache_mem_i_data[15]
+ dcache_mem_i_data[1] dcache_mem_i_data[2] dcache_mem_i_data[3] dcache_mem_i_data[4]
+ dcache_mem_i_data[5] dcache_mem_i_data[6] dcache_mem_i_data[7] dcache_mem_i_data[8]
+ dcache_mem_i_data[9] dcache_mem_o_data[0] dcache_mem_o_data[10] dcache_mem_o_data[11]
+ dcache_mem_o_data[12] dcache_mem_o_data[13] dcache_mem_o_data[14] dcache_mem_o_data[15]
+ dcache_mem_o_data[1] dcache_mem_o_data[2] dcache_mem_o_data[3] dcache_mem_o_data[4]
+ dcache_mem_o_data[5] dcache_mem_o_data[6] dcache_mem_o_data[7] dcache_mem_o_data[8]
+ dcache_mem_o_data[9] dcache_mem_req dcache_mem_sel[0] dcache_mem_sel[1] dcache_mem_we
+ dcache_rst dcache_wb_4_burst dcache_wb_ack dcache_wb_adr[0] dcache_wb_adr[10] dcache_wb_adr[11]
+ dcache_wb_adr[12] dcache_wb_adr[13] dcache_wb_adr[14] dcache_wb_adr[15] dcache_wb_adr[16]
+ dcache_wb_adr[17] dcache_wb_adr[18] dcache_wb_adr[19] dcache_wb_adr[1] dcache_wb_adr[20]
+ dcache_wb_adr[21] dcache_wb_adr[22] dcache_wb_adr[23] dcache_wb_adr[2] dcache_wb_adr[3]
+ dcache_wb_adr[4] dcache_wb_adr[5] dcache_wb_adr[6] dcache_wb_adr[7] dcache_wb_adr[8]
+ dcache_wb_adr[9] dcache_wb_cyc dcache_wb_err dcache_wb_i_dat[0] dcache_wb_i_dat[10]
+ dcache_wb_i_dat[11] dcache_wb_i_dat[12] dcache_wb_i_dat[13] dcache_wb_i_dat[14]
+ dcache_wb_i_dat[15] dcache_wb_i_dat[1] dcache_wb_i_dat[2] dcache_wb_i_dat[3] dcache_wb_i_dat[4]
+ dcache_wb_i_dat[5] dcache_wb_i_dat[6] dcache_wb_i_dat[7] dcache_wb_i_dat[8] dcache_wb_i_dat[9]
+ dcache_wb_o_dat[0] dcache_wb_o_dat[10] dcache_wb_o_dat[11] dcache_wb_o_dat[12] dcache_wb_o_dat[13]
+ dcache_wb_o_dat[14] dcache_wb_o_dat[15] dcache_wb_o_dat[1] dcache_wb_o_dat[2] dcache_wb_o_dat[3]
+ dcache_wb_o_dat[4] dcache_wb_o_dat[5] dcache_wb_o_dat[6] dcache_wb_o_dat[7] dcache_wb_o_dat[8]
+ dcache_wb_o_dat[9] dcache_wb_sel[0] dcache_wb_sel[1] dcache_wb_stb dcache_wb_we
+ ic0_clk ic0_mem_ack ic0_mem_addr[0] ic0_mem_addr[10] ic0_mem_addr[11] ic0_mem_addr[12]
+ ic0_mem_addr[13] ic0_mem_addr[14] ic0_mem_addr[15] ic0_mem_addr[1] ic0_mem_addr[2]
+ ic0_mem_addr[3] ic0_mem_addr[4] ic0_mem_addr[5] ic0_mem_addr[6] ic0_mem_addr[7]
+ ic0_mem_addr[8] ic0_mem_addr[9] ic0_mem_cache_flush ic0_mem_data[0] ic0_mem_data[10]
+ ic0_mem_data[11] ic0_mem_data[12] ic0_mem_data[13] ic0_mem_data[14] ic0_mem_data[15]
+ ic0_mem_data[16] ic0_mem_data[17] ic0_mem_data[18] ic0_mem_data[19] ic0_mem_data[1]
+ ic0_mem_data[20] ic0_mem_data[21] ic0_mem_data[22] ic0_mem_data[23] ic0_mem_data[24]
+ ic0_mem_data[25] ic0_mem_data[26] ic0_mem_data[27] ic0_mem_data[28] ic0_mem_data[29]
+ ic0_mem_data[2] ic0_mem_data[30] ic0_mem_data[31] ic0_mem_data[3] ic0_mem_data[4]
+ ic0_mem_data[5] ic0_mem_data[6] ic0_mem_data[7] ic0_mem_data[8] ic0_mem_data[9]
+ ic0_mem_ppl_submit ic0_mem_req ic0_rst ic0_wb_ack ic0_wb_adr[0] ic0_wb_adr[10] ic0_wb_adr[11]
+ ic0_wb_adr[12] ic0_wb_adr[13] ic0_wb_adr[14] ic0_wb_adr[15] ic0_wb_adr[1] ic0_wb_adr[2]
+ ic0_wb_adr[3] ic0_wb_adr[4] ic0_wb_adr[5] ic0_wb_adr[6] ic0_wb_adr[7] ic0_wb_adr[8]
+ ic0_wb_adr[9] ic0_wb_cyc ic0_wb_err ic0_wb_i_dat[0] ic0_wb_i_dat[10] ic0_wb_i_dat[11]
+ ic0_wb_i_dat[12] ic0_wb_i_dat[13] ic0_wb_i_dat[14] ic0_wb_i_dat[15] ic0_wb_i_dat[1]
+ ic0_wb_i_dat[2] ic0_wb_i_dat[3] ic0_wb_i_dat[4] ic0_wb_i_dat[5] ic0_wb_i_dat[6]
+ ic0_wb_i_dat[7] ic0_wb_i_dat[8] ic0_wb_i_dat[9] ic0_wb_sel[0] ic0_wb_sel[1] ic0_wb_stb
+ ic0_wb_we ic1_clk ic1_mem_ack ic1_mem_addr[0] ic1_mem_addr[10] ic1_mem_addr[11]
+ ic1_mem_addr[12] ic1_mem_addr[13] ic1_mem_addr[14] ic1_mem_addr[15] ic1_mem_addr[1]
+ ic1_mem_addr[2] ic1_mem_addr[3] ic1_mem_addr[4] ic1_mem_addr[5] ic1_mem_addr[6]
+ ic1_mem_addr[7] ic1_mem_addr[8] ic1_mem_addr[9] ic1_mem_cache_flush ic1_mem_data[0]
+ ic1_mem_data[10] ic1_mem_data[11] ic1_mem_data[12] ic1_mem_data[13] ic1_mem_data[14]
+ ic1_mem_data[15] ic1_mem_data[16] ic1_mem_data[17] ic1_mem_data[18] ic1_mem_data[19]
+ ic1_mem_data[1] ic1_mem_data[20] ic1_mem_data[21] ic1_mem_data[22] ic1_mem_data[23]
+ ic1_mem_data[24] ic1_mem_data[25] ic1_mem_data[26] ic1_mem_data[27] ic1_mem_data[28]
+ ic1_mem_data[29] ic1_mem_data[2] ic1_mem_data[30] ic1_mem_data[31] ic1_mem_data[3]
+ ic1_mem_data[4] ic1_mem_data[5] ic1_mem_data[6] ic1_mem_data[7] ic1_mem_data[8]
+ ic1_mem_data[9] ic1_mem_ppl_submit ic1_mem_req ic1_rst ic1_wb_ack ic1_wb_adr[0]
+ ic1_wb_adr[10] ic1_wb_adr[11] ic1_wb_adr[12] ic1_wb_adr[13] ic1_wb_adr[14] ic1_wb_adr[15]
+ ic1_wb_adr[1] ic1_wb_adr[2] ic1_wb_adr[3] ic1_wb_adr[4] ic1_wb_adr[5] ic1_wb_adr[6]
+ ic1_wb_adr[7] ic1_wb_adr[8] ic1_wb_adr[9] ic1_wb_cyc ic1_wb_err ic1_wb_i_dat[0]
+ ic1_wb_i_dat[10] ic1_wb_i_dat[11] ic1_wb_i_dat[12] ic1_wb_i_dat[13] ic1_wb_i_dat[14]
+ ic1_wb_i_dat[15] ic1_wb_i_dat[1] ic1_wb_i_dat[2] ic1_wb_i_dat[3] ic1_wb_i_dat[4]
+ ic1_wb_i_dat[5] ic1_wb_i_dat[6] ic1_wb_i_dat[7] ic1_wb_i_dat[8] ic1_wb_i_dat[9]
+ ic1_wb_sel[0] ic1_wb_sel[1] ic1_wb_stb ic1_wb_we inner_disable inner_embed_mode
+ inner_ext_irq inner_wb_4_burst inner_wb_8_burst inner_wb_ack inner_wb_adr[0] inner_wb_adr[10]
+ inner_wb_adr[11] inner_wb_adr[12] inner_wb_adr[13] inner_wb_adr[14] inner_wb_adr[15]
+ inner_wb_adr[16] inner_wb_adr[17] inner_wb_adr[18] inner_wb_adr[19] inner_wb_adr[1]
+ inner_wb_adr[20] inner_wb_adr[21] inner_wb_adr[22] inner_wb_adr[23] inner_wb_adr[2]
+ inner_wb_adr[3] inner_wb_adr[4] inner_wb_adr[5] inner_wb_adr[6] inner_wb_adr[7]
+ inner_wb_adr[8] inner_wb_adr[9] inner_wb_cyc inner_wb_err inner_wb_i_dat[0] inner_wb_i_dat[10]
+ inner_wb_i_dat[11] inner_wb_i_dat[12] inner_wb_i_dat[13] inner_wb_i_dat[14] inner_wb_i_dat[15]
+ inner_wb_i_dat[1] inner_wb_i_dat[2] inner_wb_i_dat[3] inner_wb_i_dat[4] inner_wb_i_dat[5]
+ inner_wb_i_dat[6] inner_wb_i_dat[7] inner_wb_i_dat[8] inner_wb_i_dat[9] inner_wb_o_dat[0]
+ inner_wb_o_dat[10] inner_wb_o_dat[11] inner_wb_o_dat[12] inner_wb_o_dat[13] inner_wb_o_dat[14]
+ inner_wb_o_dat[15] inner_wb_o_dat[1] inner_wb_o_dat[2] inner_wb_o_dat[3] inner_wb_o_dat[4]
+ inner_wb_o_dat[5] inner_wb_o_dat[6] inner_wb_o_dat[7] inner_wb_o_dat[8] inner_wb_o_dat[9]
+ inner_wb_sel[0] inner_wb_sel[1] inner_wb_stb inner_wb_we vccd1 vssd1
XFILLER_274_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_83_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4935__A _1999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5968__A1 _2805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3979__B1 _1462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6914_ clknet_leaf_79_core_clock _0175_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_242_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6845_ clknet_leaf_68_core_clock _0106_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_223_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4670__A _2089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6776_ clknet_leaf_85_core_clock _0037_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3988_ immu_0.page_table\[0\]\[2\] immu_0.page_table\[1\]\[2\] _1480_ vssd1 vssd1
+ vccd1 vccd1 _1500_ sky130_fd_sc_hd__mux2_1
XFILLER_183_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5727_ _2721_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_248_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3717__C _0929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6145__A1 _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5658_ _2666_ dmmu0.page_table\[11\]\[8\] _2671_ vssd1 vssd1 vccd1 vccd1 _2680_ sky130_fd_sc_hd__and3_1
XFILLER_163_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4609_ _2006_ _2047_ _2051_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__a21o_1
XFILLER_136_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5589_ _2370_ vssd1 vssd1 vccd1 vccd1 _2640_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3903__A0 _1414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7259_ clknet_leaf_25_core_clock _0520_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4548__C _2004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7061__CLK clknet_leaf_80_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6629__CLK clknet_leaf_56_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input127_A c1_o_mem_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4056__S _1390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__A3 _1483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4580__A _2017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input92_A c0_sr_bus_data_o[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4395__A0 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3293__S1 _0863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6136__A1 _2232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3696__C_N _1277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4698__A1 _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3924__A _1437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4960_ _2262_ immu_1.page_table\[7\]\[10\] _2258_ vssd1 vssd1 vccd1 vccd1 _2271_
+ sky130_fd_sc_hd__and3_1
XANTENNA__5289__C _2464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4622__A1 _2019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3911_ _1407_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__buf_6
XFILLER_205_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4891_ _2223_ vssd1 vssd1 vccd1 vccd1 _2224_ sky130_fd_sc_hd__buf_4
XFILLER_199_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4490__A _1958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6630_ clknet_leaf_55_core_clock _0700_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3842_ _1374_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5178__A2 _2390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4386__B1 inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6561_ clknet_leaf_49_core_clock _0631_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_220_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3773_ _1336_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_1
X_5512_ _2588_ immu_0.page_table\[3\]\[9\] _2591_ _2602_ vssd1 vssd1 vccd1 vccd1 _0163_
+ sky130_fd_sc_hd__a31o_1
XFILLER_185_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6492_ _3177_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4138__B1 _1535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5443_ net97 _2559_ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__and2_1
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3834__A _1363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput412 net412 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[0] sky130_fd_sc_hd__buf_2
XFILLER_145_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput423 net423 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[5] sky130_fd_sc_hd__buf_2
XFILLER_133_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6210__A _2891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput434 net434 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[14] sky130_fd_sc_hd__buf_2
X_5374_ _2310_ _2512_ vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__and2_1
XANTENNA__7084__CLK clknet_leaf_93_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput445 net445 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[24] sky130_fd_sc_hd__buf_2
Xoutput456 net456 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[5] sky130_fd_sc_hd__buf_2
XFILLER_99_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7113_ clknet_leaf_33_core_clock _0374_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[12\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3361__A1 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput467 net467 vssd1 vssd1 vccd1 vccd1 c1_i_mc_core_int sky130_fd_sc_hd__buf_2
Xoutput478 net478 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[3] sky130_fd_sc_hd__buf_2
X_4325_ _1363_ _1829_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__nor2_2
Xoutput489 net489 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[12] sky130_fd_sc_hd__buf_2
XFILLER_259_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7044_ clknet_leaf_4_core_clock _0305_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[3\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_4256_ immu_1.page_table\[8\]\[8\] immu_1.page_table\[9\]\[8\] _1524_ vssd1 vssd1
+ vccd1 vccd1 _1762_ sky130_fd_sc_hd__mux2_1
XFILLER_274_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3207_ _0818_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__4665__A _2072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4187_ _1447_ _1693_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__or2_1
XFILLER_227_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6921__CLK clknet_leaf_57_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4613__A1 _2010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5169__A2 _2390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6828_ clknet_leaf_73_core_clock _0089_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6366__A1 _3101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6759_ clknet_leaf_93_core_clock _0020_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[10\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6118__A1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3744__A _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5662__C _2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3352__A1 _0943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input244_A dcache_wb_adr[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6357__A1 _3085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5580__A2 _2632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3654__A _0901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6030__A _2879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output630_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4110_ immu_1.page_table\[8\]\[5\] immu_1.page_table\[9\]\[5\] immu_1.page_table\[10\]\[5\]
+ immu_1.page_table\[11\]\[5\] _1437_ net367 vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__mux4_2
X_5090_ _2300_ vssd1 vssd1 vccd1 vccd1 _2347_ sky130_fd_sc_hd__clkbuf_4
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4041_ _1537_ _1541_ _1542_ _1551_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__o31a_2
XFILLER_284_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4485__A _1963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4843__A1 _1981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5992_ _1968_ _2045_ vssd1 vssd1 vccd1 vccd1 _2880_ sky130_fd_sc_hd__nor2_2
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4943_ _2105_ vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__6348__A1 _3085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4874_ _2204_ immu_1.page_table\[3\]\[10\] _2196_ vssd1 vssd1 vccd1 vccd1 _2209_
+ sky130_fd_sc_hd__and3_1
XANTENNA__6205__A _2801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4651__C _2068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4359__B1 _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6613_ clknet_leaf_54_core_clock _0683_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[5\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3825_ _1365_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_1
XFILLER_192_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6544_ clknet_leaf_50_core_clock _0614_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3756_ net148 net43 _1322_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__mux2_2
XFILLER_118_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6475_ _1985_ _3157_ _3168_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__a21o_1
XFILLER_161_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3687_ dmmu1.page_table\[0\]\[11\] dmmu1.page_table\[1\]\[11\] _0856_ vssd1 vssd1
+ vccd1 vccd1 _1269_ sky130_fd_sc_hd__mux2_1
XFILLER_118_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5426_ _2546_ immu_0.page_table\[6\]\[7\] _2541_ _2551_ vssd1 vssd1 vccd1 vccd1 _0128_
+ sky130_fd_sc_hd__a31o_1
XFILLER_145_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5357_ _2503_ immu_0.page_table\[8\]\[0\] _2510_ _2511_ vssd1 vssd1 vccd1 vccd1 _0099_
+ sky130_fd_sc_hd__a31o_1
XFILLER_58_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4308_ _1584_ _1812_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__or2_1
XFILLER_141_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5288_ _2240_ _2462_ _2471_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__a21o_1
XFILLER_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5087__A1 _2332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7027_ clknet_leaf_84_core_clock _0288_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[13\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4239_ immu_0.page_table\[10\]\[8\] immu_0.page_table\[11\]\[8\] _1409_ vssd1 vssd1
+ vccd1 vccd1 _1745_ sky130_fd_sc_hd__mux2_1
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_2_0_core_clock_A clknet_1_1_1_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4047__C1 _1451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4334__S _1408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6115__A _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4561__C _2004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6817__CLK clknet_leaf_59_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input194_A c1_sr_bus_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3573__A1 _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input361_A ic1_mem_data[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3193__B _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input55_A c0_o_mem_sel[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3628__A2 _1204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4736__C _2123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6009__B _2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5848__B _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3487__S1 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6025__A _2784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output678_A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5002__A1 _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3610_ _0838_ _1193_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__nand2_1
XFILLER_266_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4590_ _2014_ _2030_ _2039_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__a21o_1
XANTENNA__5553__A2 _2623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3564__A1 _0868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3541_ _1123_ _1124_ _1125_ _0879_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__a31oi_1
XFILLER_143_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6260_ _2791_ _3040_ vssd1 vssd1 vccd1 vccd1 _3043_ sky130_fd_sc_hd__and2_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3472_ dmmu1.page_table\[0\]\[6\] dmmu1.page_table\[1\]\[6\] dmmu1.page_table\[2\]\[6\]
+ dmmu1.page_table\[3\]\[6\] _0858_ _0861_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__mux4_1
X_5211_ _2416_ dmmu0.page_table\[8\]\[8\] _2411_ vssd1 vssd1 vccd1 vccd1 _2421_ sky130_fd_sc_hd__and3_1
X_6191_ _1968_ _2255_ vssd1 vssd1 vccd1 vccd1 _3001_ sky130_fd_sc_hd__nor2_1
XFILLER_130_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5142_ _2371_ dmmu0.page_table\[10\]\[6\] _2373_ vssd1 vssd1 vccd1 vccd1 _2380_ sky130_fd_sc_hd__and3_1
XFILLER_269_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7122__CLK clknet_leaf_34_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5073_ _1930_ _2334_ vssd1 vssd1 vccd1 vccd1 _2338_ sky130_fd_sc_hd__nor2_4
XFILLER_69_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5104__A _1933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4024_ _1416_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__buf_2
XFILLER_272_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4943__A _2105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7272__CLK clknet_leaf_26_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6033__A3 _2902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5975_ _2867_ dmmu1.page_table\[13\]\[6\] _2859_ _2869_ vssd1 vssd1 vccd1 vccd1 _0359_
+ sky130_fd_sc_hd__a31o_1
X_4926_ _2237_ dmmu0.page_table\[0\]\[10\] _2220_ vssd1 vssd1 vccd1 vccd1 _2250_ sky130_fd_sc_hd__and3_1
XFILLER_240_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4857_ _2182_ immu_1.page_table\[3\]\[2\] _2197_ vssd1 vssd1 vccd1 vccd1 _2200_ sky130_fd_sc_hd__and3_1
XFILLER_220_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3993__S _1472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5774__A _2747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3808_ _1355_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_1
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4788_ _2150_ immu_1.page_table\[4\]\[4\] _2157_ vssd1 vssd1 vccd1 vccd1 _2162_ sky130_fd_sc_hd__and3_1
X_6527_ clknet_leaf_42_core_clock _0597_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3739_ net134 net29 _0847_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__mux2_1
XFILLER_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3294__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6458_ _2971_ immu_1.page_table\[8\]\[0\] _3159_ vssd1 vssd1 vccd1 vccd1 _3160_ sky130_fd_sc_hd__and3_1
XFILLER_256_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5409_ _1925_ _2540_ vssd1 vssd1 vccd1 vccd1 _2542_ sky130_fd_sc_hd__nor2_1
XFILLER_106_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6389_ net201 _3118_ vssd1 vssd1 vccd1 vccd1 _3120_ sky130_fd_sc_hd__and2_1
XFILLER_161_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5014__A _2300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4853__A _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4044__B_N _1448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6024__A3 _2877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input207_A c1_sr_bus_data_o[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5232__A1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5783__A2 _2748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_37_core_clock_A clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_169_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5299__A1 _2251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7145__CLK clknet_leaf_33_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7404__A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3932__A net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4510__A3 _1964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4239__S _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7295__CLK clknet_leaf_44_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6263__A3 _3038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5471__A1 _2576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5859__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3482__B1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5760_ _2239_ _2730_ _2740_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__a21o_1
XFILLER_201_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4711_ _2106_ immu_1.page_table\[9\]\[8\] _2103_ vssd1 vssd1 vccd1 vccd1 _2114_ sky130_fd_sc_hd__and3_1
XFILLER_194_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _2699_ vssd1 vssd1 vccd1 vccd1 _2700_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5594__A _2640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7430_ net391 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_1
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4642_ _1897_ vssd1 vssd1 vccd1 vccd1 _2072_ sky130_fd_sc_hd__buf_2
XANTENNA__3826__B net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3537__A1 _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7361_ net284 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_2
X_4573_ _1960_ _2027_ vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__or2_2
XFILLER_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3318__S _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6312_ _3069_ dmmu1.page_table\[4\]\[10\] _3057_ _3072_ vssd1 vssd1 vccd1 vccd1 _0493_
+ sky130_fd_sc_hd__a31o_1
X_3524_ _1105_ _1106_ _1108_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__nor3_1
X_7292_ clknet_leaf_43_core_clock _0553_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6243_ _3026_ dmmu1.page_table\[6\]\[8\] _3019_ _3031_ vssd1 vssd1 vccd1 vccd1 _0465_
+ sky130_fd_sc_hd__a31o_1
XFILLER_170_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3455_ _0909_ _1042_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__or2_1
XANTENNA__3842__A _1374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3396__S0 _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6174_ _2977_ dmmu1.page_table\[8\]\[6\] _2981_ _2990_ vssd1 vssd1 vccd1 vccd1 _0437_
+ sky130_fd_sc_hd__a31o_1
XFILLER_69_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3386_ _0963_ _0967_ _0972_ _0976_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__o22a_2
XANTENNA__6512__CLK clknet_leaf_58_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5125_ _2368_ vssd1 vssd1 vccd1 vccd1 _2369_ sky130_fd_sc_hd__buf_4
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5056_ _2316_ immu_0.page_table\[14\]\[5\] _2320_ _2327_ vssd1 vssd1 vccd1 vccd1
+ _0791_ sky130_fd_sc_hd__a31o_1
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3988__S _1480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5769__A _2736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4007_ _1448_ immu_1.page_table\[10\]\[2\] _1454_ vssd1 vssd1 vccd1 vccd1 _1519_
+ sky130_fd_sc_hd__o21a_1
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6662__CLK clknet_leaf_80_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6006__A3 _2878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5214__A1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5958_ _2858_ vssd1 vssd1 vccd1 vccd1 _2859_ sky130_fd_sc_hd__buf_4
XFILLER_197_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7018__CLK clknet_leaf_4_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4909_ _2237_ dmmu0.page_table\[0\]\[5\] _2221_ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__and3_1
XANTENNA__4973__B1 _2277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5889_ _2819_ dmmu0.page_table\[6\]\[4\] _2814_ vssd1 vssd1 vccd1 vccd1 _2820_ sky130_fd_sc_hd__and3_1
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7168__CLK clknet_leaf_4_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5009__A _1922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4848__A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3387__S0 _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input157_A c1_o_mem_high_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput301 ic0_mem_data[31] vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_1
Xinput312 ic0_wb_adr[12] vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_6
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput323 ic0_wb_adr[8] vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_2
Xinput334 ic1_mem_data[12] vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_2
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput345 ic1_mem_data[22] vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_2
XFILLER_248_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput356 ic1_mem_data[3] vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_2
XFILLER_263_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput367 ic1_wb_adr[13] vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_4
XANTENNA__6245__A3 _3019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input324_A ic0_wb_adr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput378 ic1_wb_adr[9] vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_2
Xinput389 inner_wb_i_dat[0] vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_16
XFILLER_263_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input18_A c0_o_mem_addr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5398__B _2527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_34_core_clock clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_189_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3199__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5756__A2 _2730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3311__S0 _0900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4192__A1 _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6535__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output543_A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4758__A _2134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3240_ net125 net20 _0840_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__mux2_1
XFILLER_112_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_73_core_clock clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__6685__CLK clknet_leaf_57_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5444__A1 _2562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5589__A _2370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4493__A _1967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6930_ clknet_leaf_77_core_clock _0191_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3550__S0 _0897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6861_ clknet_leaf_70_core_clock _0122_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5101__B _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5812_ _2223_ _2767_ _2771_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__a21o_1
XFILLER_179_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6792_ clknet_leaf_80_core_clock _0053_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5747__A2 _2730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5743_ _2729_ vssd1 vssd1 vccd1 vccd1 _2730_ sky130_fd_sc_hd__clkbuf_4
XFILLER_210_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5755__C _2732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5674_ _2210_ immu_0.high_addr_off\[0\] _2690_ vssd1 vssd1 vccd1 vccd1 _2691_ sky130_fd_sc_hd__mux2_1
XFILLER_175_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3556__B _1140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7413_ net354 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_1
X_4625_ _2054_ immu_1.page_table\[12\]\[9\] _2049_ vssd1 vssd1 vccd1 vccd1 _2060_
+ sky130_fd_sc_hd__and3_1
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7344_ net407 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4556_ _1981_ vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__buf_6
XFILLER_190_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3507_ _1089_ _1090_ _1092_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__a21oi_1
X_7275_ clknet_leaf_23_core_clock _0536_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4487_ _1965_ _1963_ vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__nor2_1
XFILLER_1_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3369__S0 _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6226_ _3010_ dmmu1.page_table\[6\]\[0\] _3019_ _3022_ vssd1 vssd1 vccd1 vccd1 _0457_
+ sky130_fd_sc_hd__a31o_1
XFILLER_103_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3438_ _0881_ _1021_ _1025_ _0887_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__a211o_1
XANTENNA__3493__A1_N _1065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6157_ _2979_ vssd1 vssd1 vccd1 vccd1 _2980_ sky130_fd_sc_hd__clkbuf_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3369_ dmmu1.page_table\[4\]\[2\] dmmu1.page_table\[5\]\[2\] dmmu1.page_table\[6\]\[2\]
+ dmmu1.page_table\[7\]\[2\] _0892_ _0864_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__mux4_1
XFILLER_97_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5108_ _1937_ _2355_ vssd1 vssd1 vccd1 vccd1 _2359_ sky130_fd_sc_hd__and2_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6088_ _2932_ dmmu1.page_table\[10\]\[11\] _2921_ _2938_ vssd1 vssd1 vccd1 vccd1
+ _0403_ sky130_fd_sc_hd__a31o_1
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5499__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5039_ _2300_ vssd1 vssd1 vccd1 vccd1 _2316_ sky130_fd_sc_hd__clkbuf_4
XFILLER_272_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6107__B _2944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4097__S1 _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3747__A _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6123__A _2216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6558__CLK clknet_leaf_50_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input274_A dcache_wb_stb vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4174__B2 _1681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4578__A _2017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput120 c1_o_mem_addr[11] vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_4
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3685__B1 _0854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput131 c1_o_mem_addr[7] vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_2
XFILLER_88_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput142 c1_o_mem_data[2] vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_2
XFILLER_248_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput153 c1_o_mem_high_addr[3] vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput164 c1_o_req_addr[0] vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_2
Xinput175 c1_o_req_addr[5] vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_1
XFILLER_263_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput186 c1_sr_bus_addr[14] vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5426__A1 _2546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput197 c1_sr_bus_data_o[0] vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_4
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5202__A _2370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5872__A _1991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4410_ net212 _0835_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__and2_1
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5390_ _2517_ immu_0.page_table\[7\]\[3\] _2525_ _2530_ vssd1 vssd1 vccd1 vccd1 _0113_
+ sky130_fd_sc_hd__a31o_1
Xoutput605 net605 vssd1 vssd1 vccd1 vccd1 ic0_rst sky130_fd_sc_hd__buf_2
Xoutput616 net616 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[2] sky130_fd_sc_hd__buf_2
Xoutput627 net627 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[11] sky130_fd_sc_hd__buf_2
XFILLER_160_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput638 net638 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[7] sky130_fd_sc_hd__buf_2
X_4341_ immu_0.page_table\[6\]\[10\] immu_0.page_table\[7\]\[10\] _1425_ vssd1 vssd1
+ vccd1 vccd1 _1845_ sky130_fd_sc_hd__mux2_1
Xoutput649 net649 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[11] sky130_fd_sc_hd__buf_2
XFILLER_207_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7060_ clknet_leaf_79_core_clock _0321_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4272_ _1581_ _1775_ _1777_ _1451_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__o211a_1
XFILLER_98_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6011_ net208 vssd1 vssd1 vccd1 vccd1 _2891_ sky130_fd_sc_hd__buf_2
XANTENNA__5665__A1 _2249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3223_ _0832_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_1
XFILLER_67_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6209__A3 _3000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4935__B _2255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6208__A _2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6090__A1 _2932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5112__A _1942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3979__A1 _1457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6913_ clknet_leaf_79_core_clock _0174_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_6844_ clknet_leaf_68_core_clock _0105_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6700__CLK clknet_leaf_42_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3987_ _1499_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_1
X_6775_ clknet_leaf_81_core_clock _0036_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5726_ immu_1.high_addr_off\[0\] _1995_ _2720_ vssd1 vssd1 vccd1 vccd1 _2721_ sky130_fd_sc_hd__mux2_1
X_5657_ _2243_ _2669_ _2679_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__a21o_1
XANTENNA__6145__A2 _2960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5782__A _2749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6850__CLK clknet_leaf_70_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4608_ _2038_ immu_1.page_table\[12\]\[1\] _2049_ vssd1 vssd1 vccd1 vccd1 _2051_
+ sky130_fd_sc_hd__and3_1
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5588_ _2233_ _2632_ _2639_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__a21o_1
XFILLER_2_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4539_ _1910_ immu_1.page_table\[14\]\[0\] _2004_ vssd1 vssd1 vccd1 vccd1 _2005_
+ sky130_fd_sc_hd__and3_1
XANTENNA__4398__A _1896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7206__CLK clknet_leaf_27_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7258_ clknet_leaf_25_core_clock _0519_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6209_ _3010_ dmmu1.page_table\[7\]\[7\] _3000_ _3011_ vssd1 vssd1 vccd1 vccd1 _0451_
+ sky130_fd_sc_hd__a31o_1
XFILLER_89_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7189_ clknet_leaf_14_core_clock _0450_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5120__A3 _2353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7502__A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4564__C _2004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5022__A _1937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3514__S0 _0896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4861__A _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4395__A1 _1894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input391_A inner_wb_i_dat[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input85_A c0_sr_bus_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6136__A2 _2960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5692__A _2443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4698__A2 _2101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6300__B _3060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4101__A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5647__A1 _2227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5111__A3 _2353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3940__A net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7412__A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6028__A _1968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_264_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6072__A1 _2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6723__CLK clknet_leaf_63_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4622__A2 _2047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4771__A _2150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3910_ _1423_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4890_ net96 vssd1 vssd1 vccd1 vccd1 _2223_ sky130_fd_sc_hd__buf_8
XFILLER_17_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3841_ _1373_ net271 vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__and2_4
XFILLER_149_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6873__CLK clknet_leaf_70_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4386__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6560_ clknet_leaf_49_core_clock _0630_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3772_ net160 net55 _0839_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__mux2_1
XANTENNA__3594__C1 _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5511_ net104 _2593_ vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__and2_1
X_6491_ dmmu1.long_off_reg\[4\] _1977_ _3172_ vssd1 vssd1 vccd1 vccd1 _3177_ sky130_fd_sc_hd__mux2_1
XANTENNA__4138__A1 _1570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5442_ _2561_ vssd1 vssd1 vccd1 vccd1 _2562_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__7229__CLK clknet_leaf_22_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3834__B net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput413 net413 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[10] sky130_fd_sc_hd__buf_2
X_5373_ _2517_ immu_0.page_table\[8\]\[7\] _2510_ _2520_ vssd1 vssd1 vccd1 vccd1 _0106_
+ sky130_fd_sc_hd__a31o_1
Xoutput424 net424 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[6] sky130_fd_sc_hd__buf_2
XFILLER_99_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6210__B _3002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput435 net435 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[15] sky130_fd_sc_hd__buf_2
Xoutput446 net446 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[25] sky130_fd_sc_hd__buf_2
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4649__C _2068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput457 net457 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[6] sky130_fd_sc_hd__buf_2
X_7112_ clknet_leaf_32_core_clock _0373_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_4324_ net107 _1810_ _1828_ _1441_ _0813_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__a221oi_1
Xoutput468 net468 vssd1 vssd1 vccd1 vccd1 c1_i_mem_ack sky130_fd_sc_hd__buf_2
XANTENNA__4011__A _1447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput479 net479 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[4] sky130_fd_sc_hd__buf_2
XFILLER_141_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7043_ clknet_leaf_17_core_clock _0304_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[3\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_4255_ _1756_ _1759_ _1760_ _1440_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__a211o_1
XANTENNA__4946__A _2262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3850__A _1378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3206_ _0823_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_1
XFILLER_234_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4186_ immu_1.page_table\[6\]\[7\] immu_1.page_table\[7\]\[7\] _1443_ vssd1 vssd1
+ vccd1 vccd1 _1693_ sky130_fd_sc_hd__mux2_1
XFILLER_255_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4613__A2 _2047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5810__A1 _2210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5777__A _2750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6827_ clknet_leaf_68_core_clock _0088_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6758_ clknet_leaf_89_core_clock _0019_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[10\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_259_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5709_ _2709_ dmmu0.page_table\[2\]\[7\] _2702_ vssd1 vssd1 vccd1 vccd1 _2711_ sky130_fd_sc_hd__and3_1
XFILLER_148_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6689_ clknet_leaf_39_core_clock _0759_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3888__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3236__S _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input237_A dcache_wb_adr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6054__A1 _2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input404_A inner_wb_i_dat[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4591__A _2038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6896__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4368__A1 _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7407__A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6311__A _2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3654__B _1235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6030__B _2904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3879__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output456_A net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4540__A1 _1996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4766__A _2134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6293__A1 _3053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4040_ _1410_ _1546_ _1550_ net315 vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_44_core_clock_A clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_256_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4843__A2 _2189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6045__A1 _2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4056__A0 _1552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5991_ net197 vssd1 vssd1 vccd1 vccd1 _2879_ sky130_fd_sc_hd__buf_2
XANTENNA__5399__A3 _2525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4942_ _1967_ _2257_ _2261_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__a21o_1
XFILLER_220_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4873_ _1987_ _2195_ _2208_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__a21o_1
XANTENNA__6205__B _3002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4359__A1 _1523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6612_ clknet_leaf_54_core_clock _0682_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[5\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3824_ _1363_ net263 vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__and2_1
XANTENNA__5556__B1 _2625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7051__CLK clknet_leaf_36_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6543_ clknet_leaf_50_core_clock _0613_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3755_ _1327_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_2
XFILLER_229_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6619__CLK clknet_leaf_53_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3845__A _1373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5763__C _2732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6474_ _2190_ immu_1.page_table\[8\]\[8\] _3159_ vssd1 vssd1 vccd1 vccd1 _3168_ sky130_fd_sc_hd__and3_1
X_3686_ _1261_ _1263_ _1265_ _1267_ net123 vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__o221a_2
XFILLER_173_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5425_ net102 _2543_ vssd1 vssd1 vccd1 vccd1 _2551_ sky130_fd_sc_hd__and2_1
XFILLER_160_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5323__A3 _2480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3283__C net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5356_ _1926_ _2509_ vssd1 vssd1 vccd1 vccd1 _2511_ sky130_fd_sc_hd__nor2_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4307_ immu_1.page_table\[14\]\[9\] immu_1.page_table\[15\]\[9\] _1453_ vssd1 vssd1
+ vccd1 vccd1 _1812_ sky130_fd_sc_hd__mux2_1
XANTENNA__4676__A _2089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5287_ _2458_ dmmu0.page_table\[14\]\[6\] _2464_ vssd1 vssd1 vccd1 vccd1 _2471_ sky130_fd_sc_hd__and3_1
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6284__A1 _3053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7026_ clknet_leaf_82_core_clock _0287_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_4238_ _1570_ _1741_ _1743_ _1535_ vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__o211a_1
XFILLER_101_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4169_ net112 immu_1.high_addr_off\[2\] vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__nand2_1
XFILLER_228_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5003__C _2282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4598__A1 _2023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5300__A _2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6115__B _2944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3755__A _1327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6131__A _2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input187_A c1_sr_bus_addr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5314__A3 _2480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input354_A ic1_mem_data[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4522__A1 _1976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3193__C net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3956__S0 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input48_A c0_o_mem_high_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4586__A _2017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6275__A1 _3042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4038__B1 _1416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6306__A _2931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4752__C _2140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7074__CLK clknet_leaf_79_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6025__B _2064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5002__A2 _2280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5223__A_N _2367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4260__S _1524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5583__C _2634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3540_ _1090_ _1092_ _1089_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__a21bo_1
XANTENNA__4761__A1 _2012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6911__CLK clknet_leaf_76_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3471_ dmmu1.page_table\[4\]\[6\] dmmu1.page_table\[5\]\[6\] dmmu1.page_table\[6\]\[6\]
+ dmmu1.page_table\[7\]\[6\] _0858_ _0861_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__mux4_1
XFILLER_142_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5305__A3 _2480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5880__A _2777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5210_ _2243_ _2409_ _2420_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__a21o_1
XFILLER_142_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4513__A1 _1976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6190_ _2999_ vssd1 vssd1 vccd1 vccd1 _3000_ sky130_fd_sc_hd__buf_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5141_ _2236_ _2369_ _2379_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a21o_1
XFILLER_130_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4496__A _1972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5072_ _2332_ immu_0.page_table\[12\]\[0\] _2336_ _2337_ vssd1 vssd1 vccd1 vccd1
+ _0797_ sky130_fd_sc_hd__a31o_1
XFILLER_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4023_ _1534_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5104__B _2355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6216__A _1991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5974_ _2801_ _2861_ vssd1 vssd1 vccd1 vccd1 _2869_ sky130_fd_sc_hd__and2_1
XFILLER_225_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4925_ _1950_ vssd1 vssd1 vccd1 vccd1 _2249_ sky130_fd_sc_hd__buf_4
X_4856_ _1967_ _2195_ _2199_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__a21o_1
XFILLER_178_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3807_ net217 _1348_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__and2_1
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4787_ _2010_ _2155_ _2161_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__a21o_1
X_6526_ clknet_leaf_30_core_clock _0596_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[14\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3738_ _1318_ vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_4
XFILLER_109_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6591__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6457_ _3158_ vssd1 vssd1 vccd1 vccd1 _3159_ sky130_fd_sc_hd__buf_2
XFILLER_69_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3669_ net51 dmmu0.long_off_reg\[6\] vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__and2_1
XFILLER_106_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5790__A _2749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4504__A1 _1976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5408_ _2540_ vssd1 vssd1 vccd1 vccd1 _2541_ sky130_fd_sc_hd__clkbuf_4
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6388_ _3112_ dmmu1.page_table\[1\]\[0\] _3116_ _3119_ vssd1 vssd1 vccd1 vccd1 _0522_
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5339_ _1937_ _2497_ vssd1 vssd1 vccd1 vccd1 _2501_ sky130_fd_sc_hd__and2_1
XFILLER_114_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7009_ clknet_leaf_78_core_clock _0270_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7097__CLK clknet_leaf_36_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_core_clock clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4345__S _1425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5668__C _2670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5030__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5232__A2 _2430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input102_A c0_sr_bus_data_o[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5965__A _2793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6934__CLK clknet_leaf_75_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5535__A3 _2607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4743__A1 _2023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5205__A _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_63_core_clock clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4259__B1 _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7420__A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6036__A _2795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6420__A1 _3128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4710_ _2019_ _2101_ _2113_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__a21o_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _2217_ _2605_ vssd1 vssd1 vccd1 vccd1 _2699_ sky130_fd_sc_hd__nor2_1
X_4641_ _2008_ _2066_ _2071_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__a21o_1
X_4572_ net188 net181 vssd1 vssd1 vccd1 vccd1 _2027_ sky130_fd_sc_hd__or2b_1
X_7360_ net283 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__buf_2
XFILLER_128_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6311_ _2895_ _3059_ vssd1 vssd1 vccd1 vccd1 _3072_ sky130_fd_sc_hd__and2_1
X_3523_ _1105_ _1106_ _1108_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__o21a_1
X_7291_ clknet_leaf_44_core_clock _0552_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6487__A1 _1972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6242_ _2891_ _3021_ vssd1 vssd1 vccd1 vccd1 _3031_ sky130_fd_sc_hd__and2_1
X_3454_ dmmu0.page_table\[2\]\[5\] dmmu0.page_table\[3\]\[5\] _0910_ vssd1 vssd1 vccd1
+ vccd1 _1042_ sky130_fd_sc_hd__mux2_1
XFILLER_143_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6173_ _2801_ _2983_ vssd1 vssd1 vccd1 vccd1 _2990_ sky130_fd_sc_hd__and2_1
X_3385_ _0918_ _0929_ _0975_ _0835_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__a31o_1
XANTENNA__3396__S1 _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6239__A1 _3026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5124_ _2217_ _2367_ vssd1 vssd1 vccd1 vccd1 _2368_ sky130_fd_sc_hd__nor2_1
XFILLER_97_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5055_ _1940_ _2322_ vssd1 vssd1 vccd1 vccd1 _2327_ sky130_fd_sc_hd__and2_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4954__A _2262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6807__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4006_ immu_1.page_table\[11\]\[2\] _1448_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__or2b_1
XFILLER_242_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6411__A1 _3128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5214__A2 _2409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6957__CLK clknet_leaf_81_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5957_ _2857_ vssd1 vssd1 vccd1 vccd1 _2858_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_201_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4908_ _2105_ vssd1 vssd1 vccd1 vccd1 _2237_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__4973__A1 _1979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5888_ _2681_ vssd1 vssd1 vccd1 vccd1 _2819_ sky130_fd_sc_hd__buf_2
X_4839_ _1972_ _2189_ _2192_ immu_1.page_table\[1\]\[2\] vssd1 vssd1 vccd1 vccd1 _0709_
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4725__A1 _1996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5009__B _2296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6509_ clknet_leaf_59_core_clock _0579_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7489_ net109 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_1
XANTENNA__7505__A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4848__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3387__S1 _0864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3244__S _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4567__C _2004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput302 ic0_mem_data[3] vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_1
Xinput313 ic0_wb_adr[13] vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_4
XFILLER_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput324 ic0_wb_adr[9] vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput335 ic1_mem_data[13] vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_2
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput346 ic1_mem_data[23] vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_2
Xinput357 ic1_mem_data[4] vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_2
XFILLER_152_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput368 ic1_wb_adr[14] vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_2
Xinput379 ic1_wb_cyc vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input317_A ic0_wb_adr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3464__A1 _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4075__S _1438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6402__A1 _3112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3199__B _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3311__S1 _0902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3927__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5508__A3 _2591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7112__CLK clknet_leaf_32_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4716__A1 _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6469__A1 _1979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3943__A net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7262__CLK clknet_leaf_25_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5141__A1 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output536_A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4493__B _1970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5995__A3 _2878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6860_ clknet_leaf_71_core_clock _0121_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3550__S1 _0902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5811_ _2762_ dmmu0.page_table\[3\]\[1\] _2769_ vssd1 vssd1 vccd1 vccd1 _2771_ sky130_fd_sc_hd__and3_1
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6791_ clknet_leaf_80_core_clock _0052_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5742_ _2216_ _2572_ vssd1 vssd1 vccd1 vccd1 _2729_ sky130_fd_sc_hd__nor2_2
XANTENNA__4955__A1 _1983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5673_ _2689_ vssd1 vssd1 vccd1 vccd1 _2690_ sky130_fd_sc_hd__buf_4
XFILLER_148_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7412_ net352 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_1
X_4624_ _2021_ _2047_ _2059_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__a21o_1
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6172__A3 _2981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7343_ net386 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_4
XFILLER_190_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4555_ _2014_ _2002_ _2015_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__a21o_1
XFILLER_116_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3853__A _1373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3506_ net150 dmmu1.long_off_reg\[0\] _1066_ _1091_ vssd1 vssd1 vccd1 vccd1 _1092_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__5771__C _2731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7274_ clknet_leaf_20_core_clock _0535_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4486_ net197 vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__inv_2
XFILLER_116_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6225_ _2879_ _3021_ vssd1 vssd1 vccd1 vccd1 _3022_ sky130_fd_sc_hd__and2_1
XFILLER_249_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3437_ _0869_ _1022_ _1024_ _0855_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__o211a_1
XANTENNA__3369__S1 _0864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6156_ _2919_ _2978_ vssd1 vssd1 vccd1 vccd1 _2979_ sky130_fd_sc_hd__or2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _0819_ _0944_ _0956_ _0959_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__a22o_2
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3694__A1 _0868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3999__S _1472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _2347_ immu_0.page_table\[13\]\[3\] _2353_ _2358_ vssd1 vssd1 vccd1 vccd1
+ _0002_ sky130_fd_sc_hd__a31o_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4684__A _2089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6087_ _1991_ _2923_ vssd1 vssd1 vccd1 vccd1 _2938_ sky130_fd_sc_hd__and2_1
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3299_ _0891_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__buf_6
XFILLER_181_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5499__B _2593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5038_ _2301_ immu_0.page_table\[15\]\[10\] _2297_ _2315_ vssd1 vssd1 vccd1 vccd1
+ _0785_ sky130_fd_sc_hd__a31o_1
XFILLER_122_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5199__A1 _2227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6989_ clknet_leaf_7_core_clock _0250_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7135__CLK clknet_leaf_34_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6123__B _2621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7285__CLK clknet_leaf_26_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5371__A1 _2517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4174__A2 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4859__A _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3763__A _1331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input267_A dcache_wb_o_dat[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3685__A1 _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput110 c1_o_instr_long_addr[0] vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_2
XFILLER_248_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput121 c1_o_mem_addr[12] vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_4
XFILLER_264_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput132 c1_o_mem_addr[8] vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_2
XANTENNA_input30_A c0_o_mem_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput143 c1_o_mem_data[3] vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_2
Xinput154 c1_o_mem_high_addr[4] vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_1
XFILLER_264_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput165 c1_o_req_addr[10] vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_1
Xinput176 c1_o_req_addr[6] vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput187 c1_sr_bus_addr[15] vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_49_core_clock_A clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput198 c1_sr_bus_data_o[10] vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_4
XANTENNA__3437__A1 _0869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5977__A3 _2859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4760__C _2140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output486_A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5362__A1 _2503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput606 net606 vssd1 vssd1 vccd1 vccd1 ic0_wb_ack sky130_fd_sc_hd__buf_2
XFILLER_160_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6652__CLK clknet_leaf_38_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput617 net617 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[3] sky130_fd_sc_hd__buf_2
XFILLER_125_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput628 net628 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[12] sky130_fd_sc_hd__buf_2
X_4340_ _1837_ _1839_ _1841_ _1843_ _1413_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__o221a_1
XFILLER_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput639 net639 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[8] sky130_fd_sc_hd__buf_2
XFILLER_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4271_ _1447_ _1776_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__or2_1
XFILLER_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6010_ _2884_ dmmu1.page_table\[12\]\[7\] _2878_ _2890_ vssd1 vssd1 vccd1 vccd1 _0373_
+ sky130_fd_sc_hd__a31o_1
X_3222_ net216 _0824_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__and2_1
XANTENNA__7008__CLK clknet_leaf_79_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6208__B _3002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5968__A3 _2859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5112__B _2355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6912_ clknet_leaf_72_core_clock _0173_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__7158__CLK clknet_leaf_12_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6843_ clknet_leaf_68_core_clock _0104_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3848__A _1377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6224__A _3020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6774_ clknet_leaf_91_core_clock _0035_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[9\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4670__C _2086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3986_ net235 _1498_ _0811_ vssd1 vssd1 vccd1 vccd1 _1499_ sky130_fd_sc_hd__mux2_4
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5725_ _1997_ _2719_ vssd1 vssd1 vccd1 vccd1 _2720_ sky130_fd_sc_hd__nor2_8
XFILLER_50_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_51_core_clock_A clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5656_ _2666_ dmmu0.page_table\[11\]\[7\] _2671_ vssd1 vssd1 vccd1 vccd1 _2679_ sky130_fd_sc_hd__and3_1
XFILLER_108_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4607_ _1996_ _2047_ _2050_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__a21o_1
XANTENNA__5353__A1 _2503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5587_ _2473_ dmmu0.page_table\[12\]\[4\] _2634_ vssd1 vssd1 vccd1 vccd1 _2639_ sky130_fd_sc_hd__and3_1
XFILLER_151_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4538_ _2003_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__clkbuf_4
XFILLER_264_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5105__A1 _2347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7257_ clknet_leaf_25_core_clock _0518_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4469_ _1939_ immu_0.page_table\[11\]\[9\] _1924_ _1949_ vssd1 vssd1 vccd1 vccd1
+ _0582_ sky130_fd_sc_hd__a31o_1
XFILLER_277_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4313__C1 _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6208_ _2803_ _3002_ vssd1 vssd1 vccd1 vccd1 _3011_ sky130_fd_sc_hd__and2_1
XFILLER_131_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7188_ clknet_leaf_14_core_clock _0449_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_258_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _2845_ dmmu0.page_table\[1\]\[6\] _2962_ vssd1 vssd1 vccd1 vccd1 _2969_ sky130_fd_sc_hd__and3_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5022__B _2302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3514__S1 _0901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4580__C _2032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6675__CLK clknet_leaf_56_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input384_A inner_disable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5692__B _2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4589__A _2038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input78_A c0_sr_bus_addr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5647__A2 _2669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3658__A1 dmmu0.page_table\[9\]\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6309__A _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7300__CLK clknet_leaf_44_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5213__A _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6028__B _2064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6044__A _2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3840_ inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3269__S0 _0858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3771_ _1335_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_1
XFILLER_220_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5510_ _2588_ immu_0.page_table\[3\]\[8\] _2591_ _2601_ vssd1 vssd1 vccd1 vccd1 _0162_
+ sky130_fd_sc_hd__a31o_1
XFILLER_285_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6490_ _3176_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4138__A2 _1645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5441_ _1897_ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__buf_4
XFILLER_157_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4499__A _1974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3346__B1 _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput414 net414 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[11] sky130_fd_sc_hd__buf_2
XFILLER_160_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5372_ _1944_ _2512_ vssd1 vssd1 vccd1 vccd1 _2520_ sky130_fd_sc_hd__and2_1
Xoutput425 net425 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[7] sky130_fd_sc_hd__buf_2
XFILLER_172_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput436 net436 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[16] sky130_fd_sc_hd__buf_2
X_7111_ clknet_leaf_35_core_clock _0372_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput447 net447 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[26] sky130_fd_sc_hd__buf_2
X_4323_ _1457_ _1814_ _1818_ _1822_ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__o32a_1
Xoutput458 net458 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[7] sky130_fd_sc_hd__buf_2
XFILLER_141_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput469 net469 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[0] sky130_fd_sc_hd__buf_2
XFILLER_259_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7042_ clknet_leaf_17_core_clock _0303_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4254_ _1684_ _1757_ _1758_ _1756_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__a22oi_1
XANTENNA__4846__B1 _2192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3205_ net223 _0819_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__and2_1
XFILLER_228_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4185_ immu_1.page_table\[4\]\[7\] immu_1.page_table\[5\]\[7\] _1493_ vssd1 vssd1
+ vccd1 vccd1 _1692_ sky130_fd_sc_hd__mux2_1
XANTENNA__4665__C _2086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6548__CLK clknet_leaf_48_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4962__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3282__C1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6698__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6826_ clknet_leaf_60_core_clock _0087_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[10\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_250_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6366__A3 _3096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6757_ clknet_leaf_90_core_clock _0018_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[10\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5574__A1 _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3969_ _1479_ _1481_ _1411_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__o21ai_1
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5708_ _2240_ _2700_ _2710_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__a21o_1
XFILLER_136_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6688_ clknet_leaf_56_core_clock _0758_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5639_ _2668_ vssd1 vssd1 vccd1 vccd1 _2669_ sky130_fd_sc_hd__buf_4
XANTENNA__6401__B _3118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3337__A0 _0898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3888__A1 _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7309_ clknet_leaf_19_core_clock _0570_ vssd1 vssd1 vccd1 vccd1 dmmu1.long_off_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5732__S _2720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4837__B1 _2192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6129__A _2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5033__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input132_A c1_o_mem_addr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4872__A _2204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4065__A1 _1572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6357__A3 _3096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5565__A1 _2223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3576__B1 _0854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6311__B _3059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3879__A1 _1397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4540__A2 _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output449_A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7423__A net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4258__S _1493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5878__A _2443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4782__A _2150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5990_ _2877_ vssd1 vssd1 vccd1 vccd1 _2878_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__6840__CLK clknet_leaf_69_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4056__A1 _1566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4941_ _2237_ immu_1.page_table\[7\]\[1\] _2259_ vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__and3_1
XFILLER_212_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4872_ _2204_ immu_1.page_table\[3\]\[9\] _2197_ vssd1 vssd1 vccd1 vccd1 _2208_ sky130_fd_sc_hd__and3_1
XFILLER_60_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6611_ clknet_leaf_53_core_clock _0681_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3823_ _1364_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5556__A1 _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6542_ clknet_leaf_48_core_clock _0612_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3754_ net147 net42 _1322_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__mux2_2
XFILLER_118_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5308__A1 _2363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6473_ _1983_ _3157_ _3167_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__a21o_1
X_3685_ _0859_ _1266_ _0854_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__o21ai_1
XANTENNA__3337__S _0929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5424_ _2546_ immu_0.page_table\[6\]\[6\] _2541_ _2550_ vssd1 vssd1 vccd1 vccd1 _0127_
+ sky130_fd_sc_hd__a31o_1
XFILLER_133_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3414__S0 _0865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5355_ _2509_ vssd1 vssd1 vccd1 vccd1 _2510_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3283__D net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4306_ immu_1.page_table\[12\]\[9\] immu_1.page_table\[13\]\[9\] _1524_ vssd1 vssd1
+ vccd1 vccd1 _1811_ sky130_fd_sc_hd__mux2_1
XFILLER_245_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5286_ _2236_ _2462_ _2470_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__a21o_1
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7025_ clknet_leaf_83_core_clock _0286_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5087__A3 _2336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4237_ _1478_ _1742_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__or2_1
XFILLER_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4168_ net112 immu_1.high_addr_off\[2\] vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__nor2_1
XFILLER_255_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5788__A _2749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_core_clock clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_243_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4099_ _1479_ _1605_ _1607_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__a21o_1
XANTENNA__4047__B2 _1447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4598__A2 _2030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5795__A1 _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6809_ clknet_leaf_86_core_clock _0070_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7508__A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6412__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6131__B dmmu0.page_table\[1\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5028__A _1944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3956__S1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3771__A _1335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_core_clock clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_105_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input347_A ic1_mem_data[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6863__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5698__A _2682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4038__A1 _1419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5235__B1 _1911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7219__CLK clknet_leaf_27_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4107__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7418__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3549__B1 _0957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6322__A _2879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4761__A2 _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3470_ _0993_ _1035_ _1054_ _1057_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__o22a_4
XFILLER_170_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5710__A1 _2243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5140_ _2371_ dmmu0.page_table\[10\]\[5\] _2373_ vssd1 vssd1 vccd1 vccd1 _2379_ sky130_fd_sc_hd__and3_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4496__B _1970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5071_ _1926_ _2335_ vssd1 vssd1 vccd1 vccd1 _2337_ sky130_fd_sc_hd__nor2_1
XFILLER_84_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4022_ net236 _1533_ _0811_ vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__mux2_4
XFILLER_231_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5973_ _2867_ dmmu1.page_table\[13\]\[5\] _2859_ _2868_ vssd1 vssd1 vccd1 vccd1 _0358_
+ sky130_fd_sc_hd__a31o_1
XFILLER_252_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4924_ _2247_ _2219_ _2248_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__a21o_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5529__A1 _2603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4855_ _2182_ immu_1.page_table\[3\]\[1\] _2197_ vssd1 vssd1 vccd1 vccd1 _2199_ sky130_fd_sc_hd__and3_1
XFILLER_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3806_ _1354_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_1
XFILLER_220_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4786_ _2150_ immu_1.page_table\[4\]\[3\] _2157_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__and3_1
XANTENNA__3635__S0 _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6736__CLK clknet_leaf_66_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6525_ clknet_leaf_31_core_clock _0595_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[14\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_3737_ _1299_ _1317_ _0818_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__mux2_1
X_6456_ _2084_ _2978_ vssd1 vssd1 vccd1 vccd1 _3158_ sky130_fd_sc_hd__or2_1
X_3668_ net51 dmmu0.long_off_reg\[6\] vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__nor2_1
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5407_ _1929_ _2539_ vssd1 vssd1 vccd1 vccd1 _2540_ sky130_fd_sc_hd__or2_1
XFILLER_161_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5701__A1 _2230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6387_ net197 _3118_ vssd1 vssd1 vccd1 vccd1 _3119_ sky130_fd_sc_hd__and2_1
XANTENNA__3591__A _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6886__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3599_ dmmu0.page_table\[2\]\[9\] dmmu0.page_table\[3\]\[9\] _1169_ vssd1 vssd1 vccd1
+ vccd1 _1183_ sky130_fd_sc_hd__mux2_1
X_5338_ _2489_ immu_0.page_table\[9\]\[3\] _2495_ _2500_ vssd1 vssd1 vccd1 vccd1 _0091_
+ sky130_fd_sc_hd__a31o_1
XFILLER_272_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5269_ _2458_ dmmu0.page_table\[7\]\[12\] _2444_ vssd1 vssd1 vccd1 vccd1 _2460_ sky130_fd_sc_hd__and3_1
XFILLER_272_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7008_ clknet_leaf_79_core_clock _0269_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_263_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3530__S _0854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5311__A _1935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4853__C _2197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5768__A1 _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5965__B _2861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4361__S _1524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input297_A ic0_mem_data[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4743__A2 _2120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5940__A1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3951__B1 _1464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input60_A c0_o_req_addr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4597__A _2038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4259__A1 _1523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5471__A3 _2574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6609__CLK clknet_leaf_53_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6317__A _2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3440__S _0865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6036__B _2904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7191__CLK clknet_leaf_28_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6759__CLK clknet_leaf_93_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4640_ _2054_ immu_1.page_table\[11\]\[2\] _2068_ vssd1 vssd1 vccd1 vccd1 _2071_
+ sky130_fd_sc_hd__and3_1
XFILLER_202_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5594__C _2634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4571_ _2025_ _2001_ _2026_ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__a21o_1
XFILLER_190_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5931__A1 _1948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5891__A _2819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6310_ _3069_ dmmu1.page_table\[4\]\[9\] _3058_ _3071_ vssd1 vssd1 vccd1 vccd1 _0492_
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_56_core_clock_A clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3522_ net45 dmmu0.long_off_reg\[0\] _1077_ _1107_ vssd1 vssd1 vccd1 vccd1 _1108_
+ sky130_fd_sc_hd__a31oi_2
X_7290_ clknet_leaf_92_core_clock _0551_ vssd1 vssd1 vccd1 vccd1 mem_dcache_arb.transfer_active
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6241_ _3026_ dmmu1.page_table\[6\]\[7\] _3019_ _3030_ vssd1 vssd1 vccd1 vccd1 _0464_
+ sky130_fd_sc_hd__a31o_1
X_3453_ _0948_ _1040_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__or2_1
XFILLER_170_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6172_ _2977_ dmmu1.page_table\[8\]\[5\] _2981_ _2989_ vssd1 vssd1 vccd1 vccd1 _0436_
+ sky130_fd_sc_hd__a31o_1
X_3384_ _0973_ _0974_ _0899_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__mux2_1
XFILLER_226_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5123_ _1913_ _2317_ vssd1 vssd1 vccd1 vccd1 _2367_ sky130_fd_sc_hd__or2_4
XFILLER_69_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _2316_ immu_0.page_table\[14\]\[4\] _2320_ _2326_ vssd1 vssd1 vccd1 vccd1
+ _0790_ sky130_fd_sc_hd__a31o_1
XFILLER_238_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4005_ immu_1.page_table\[0\]\[2\] immu_1.page_table\[1\]\[2\] immu_1.page_table\[2\]\[2\]
+ immu_1.page_table\[3\]\[2\] _1453_ _1454_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__mux4_1
XFILLER_284_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6227__A _2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5769__C _2731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5956_ _2784_ _2028_ vssd1 vssd1 vccd1 vccd1 _2857_ sky130_fd_sc_hd__or2_1
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4907_ _2235_ vssd1 vssd1 vccd1 vccd1 _2236_ sky130_fd_sc_hd__buf_4
XFILLER_200_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5887_ _2229_ _2812_ _2818_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__a21o_1
XANTENNA__4973__A2 _2274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4181__S _1493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4838_ _1967_ _2189_ _2192_ immu_1.page_table\[1\]\[1\] vssd1 vssd1 vccd1 vccd1 _0708_
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4725__A2 _2120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4769_ _2021_ _2138_ _2149_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__a21o_1
XFILLER_193_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6508_ clknet_leaf_60_core_clock _0578_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_106_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7488_ net170 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_2
XFILLER_134_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6439_ net198 _3136_ vssd1 vssd1 vccd1 vccd1 _3148_ sky130_fd_sc_hd__and2_1
XFILLER_134_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5686__A0 _2239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5306__A _1930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7064__CLK clknet_leaf_10_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_core_clock clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_core_clock
+ sky130_fd_sc_hd__clkbuf_16
Xinput303 ic0_mem_data[4] vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput314 ic0_wb_adr[14] vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_2
XANTENNA__5740__S _2720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput325 ic0_wb_cyc vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_2
Xinput336 ic1_mem_data[14] vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_2
Xinput347 ic1_mem_data[24] vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__buf_2
XFILLER_75_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput358 ic1_mem_data[5] vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_2
XFILLER_152_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput369 ic1_wb_adr[15] vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_4
XFILLER_248_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4356__S _1439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6137__A _2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input212_A dcache_mem_ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5976__A _2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6166__A1 _2977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_4_0_core_clock clknet_2_2_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_125_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6469__A2 _3157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3435__S _0857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4758__C _2140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5141__A2 _2369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output431_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output529_A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7431__A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5444__A3 _2557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4652__A1 _2019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6581__CLK clknet_leaf_46_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5886__A _2777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5810_ _2210_ _2767_ _2770_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__a21o_1
XFILLER_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4790__A _2150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6790_ clknet_leaf_80_core_clock _0051_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_5741_ _2728_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4955__A2 _2257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5672_ _1917_ _2688_ vssd1 vssd1 vccd1 vccd1 _2689_ sky130_fd_sc_hd__or2_1
XFILLER_175_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7411_ net351 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_1
X_4623_ _2054_ immu_1.page_table\[12\]\[8\] _2049_ vssd1 vssd1 vccd1 vccd1 _2059_
+ sky130_fd_sc_hd__and3_1
XFILLER_148_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5904__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7342_ net384 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_1
X_4554_ _1910_ immu_1.page_table\[14\]\[5\] _2004_ vssd1 vssd1 vccd1 vccd1 _2015_
+ sky130_fd_sc_hd__and3_1
XFILLER_128_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7087__CLK clknet_leaf_93_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3505_ net151 dmmu1.long_off_reg\[1\] vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__and2_1
X_7273_ clknet_leaf_26_core_clock _0534_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_4485_ _1963_ vssd1 vssd1 vccd1 vccd1 _1964_ sky130_fd_sc_hd__clkbuf_4
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5126__A _1896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6224_ _3020_ vssd1 vssd1 vccd1 vccd1 _3021_ sky130_fd_sc_hd__clkbuf_4
XFILLER_116_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3436_ _0863_ _1023_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__or2_1
XFILLER_131_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4340__B1 _1841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6155_ net188 net181 _2062_ vssd1 vssd1 vccd1 vccd1 _2978_ sky130_fd_sc_hd__or3_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4965__A _2190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _0909_ _0958_ _0819_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__a21oi_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7341__A clknet_leaf_92_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _1935_ _2355_ vssd1 vssd1 vccd1 vccd1 _2358_ sky130_fd_sc_hd__and2_1
XFILLER_111_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6086_ _2932_ dmmu1.page_table\[10\]\[10\] _2921_ _2937_ vssd1 vssd1 vccd1 vccd1
+ _0402_ sky130_fd_sc_hd__a31o_1
XFILLER_257_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3298_ _0857_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__buf_6
XANTENNA__6924__CLK clknet_leaf_58_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5037_ _2314_ _2302_ vssd1 vssd1 vccd1 vccd1 _2315_ sky130_fd_sc_hd__and2_1
XFILLER_272_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5796__A _2749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6396__A1 _3112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5199__A2 _2409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6988_ clknet_leaf_8_core_clock _0249_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_213_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5939_ _2214_ _2688_ vssd1 vssd1 vccd1 vccd1 _2848_ sky130_fd_sc_hd__nor2_4
XFILLER_15_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3382__A1 dmmu0.page_table\[1\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3255__S _0847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4578__C _2032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5036__A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input162_A c1_o_mem_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput100 c0_sr_bus_data_o[5] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__buf_6
XFILLER_88_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput111 c1_o_instr_long_addr[1] vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_2
Xinput122 c1_o_mem_addr[13] vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_2
XFILLER_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput133 c1_o_mem_addr[9] vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_2
Xinput144 c1_o_mem_data[4] vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
XFILLER_236_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput155 c1_o_mem_high_addr[5] vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput166 c1_o_req_addr[11] vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_1
XFILLER_276_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput177 c1_o_req_addr[7] vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input23_A c0_o_mem_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5426__A3 _2541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput188 c1_sr_bus_addr[1] vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_4
XFILLER_236_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput199 c1_sr_bus_data_o[11] vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_2
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3954__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7426__A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6330__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput607 net607 vssd1 vssd1 vccd1 vccd1 ic0_wb_err sky130_fd_sc_hd__buf_2
Xoutput618 net618 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[4] sky130_fd_sc_hd__buf_2
XFILLER_172_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput629 net629 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[13] sky130_fd_sc_hd__buf_2
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4270_ immu_1.page_table\[2\]\[8\] immu_1.page_table\[3\]\[8\] _1437_ vssd1 vssd1
+ vccd1 vccd1 _1776_ sky130_fd_sc_hd__mux2_1
XFILLER_207_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6947__CLK clknet_leaf_1_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4322__B1 _1553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3221_ _0831_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4873__A1 _1987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6911_ clknet_leaf_76_core_clock _0172_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6378__A1 _3101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6842_ clknet_leaf_69_core_clock _0103_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4389__A0 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6773_ clknet_leaf_91_core_clock _0034_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[9\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3985_ _0813_ _1477_ _1483_ _1497_ vssd1 vssd1 vccd1 vccd1 _1498_ sky130_fd_sc_hd__a31o_1
XANTENNA__5050__A1 _2316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5724_ net710 _2718_ _1955_ _2272_ vssd1 vssd1 vccd1 vccd1 _2719_ sky130_fd_sc_hd__or4_4
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5655_ _2240_ _2669_ _2678_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__a21o_1
XANTENNA__3864__A _1387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4606_ _2038_ immu_1.page_table\[12\]\[0\] _2049_ vssd1 vssd1 vccd1 vccd1 _2050_
+ sky130_fd_sc_hd__and3_1
XFILLER_190_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6240__A _2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5782__C _2751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5586_ _2230_ _2632_ _2638_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__a21o_1
XANTENNA__4010__C1 _1441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4537_ _1961_ _1998_ vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__or2_1
XFILLER_190_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7256_ clknet_leaf_24_core_clock _0517_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4468_ _1948_ _1931_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__and2_1
XFILLER_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6207_ _2931_ vssd1 vssd1 vccd1 vccd1 _3010_ sky130_fd_sc_hd__buf_4
XFILLER_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3419_ _0924_ _0925_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__nor2_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4695__A _1896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7187_ clknet_leaf_28_core_clock _0448_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4399_ _1897_ vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__buf_6
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4864__A1 _1979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6138_ _2235_ _2960_ _2968_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__a21o_1
XFILLER_246_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7102__CLK clknet_leaf_30_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6069_ _2795_ _2924_ vssd1 vssd1 vccd1 vccd1 _2928_ sky130_fd_sc_hd__and2_1
XFILLER_280_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4616__A1 _2012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4077__C1 _1516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4861__C _2197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6150__A _2971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input377_A ic1_wb_adr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4001__C1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_opt_2_0_core_clock clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_opt_2_0_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_181_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_7_0_core_clock_A clknet_2_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_107_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3713__S net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6309__B _3060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4607__A1 _1996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6072__A3 _2922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5280__A1 _2227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4771__C _2140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6044__B _2904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5032__A1 _2301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3269__S1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3770_ net140 net35 _0839_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__mux2_8
XFILLER_192_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5440_ _2546_ immu_0.page_table\[5\]\[1\] _2557_ _2560_ vssd1 vssd1 vccd1 vccd1 _0133_
+ sky130_fd_sc_hd__a31o_1
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4499__B _1970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3346__A1 _0881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5371_ _2517_ immu_0.page_table\[8\]\[6\] _2510_ _2519_ vssd1 vssd1 vccd1 vccd1 _0105_
+ sky130_fd_sc_hd__a31o_1
Xoutput415 net415 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[12] sky130_fd_sc_hd__buf_2
XFILLER_126_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput426 net426 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[8] sky130_fd_sc_hd__buf_2
Xoutput437 net437 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[17] sky130_fd_sc_hd__buf_2
X_7110_ clknet_leaf_35_core_clock _0371_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4322_ _1530_ _1824_ _1826_ _1553_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__a31o_1
Xoutput448 net448 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[27] sky130_fd_sc_hd__buf_2
Xoutput459 net459 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[8] sky130_fd_sc_hd__buf_2
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7041_ clknet_leaf_17_core_clock _0302_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_4253_ _1684_ _1757_ _1758_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__and3_1
XANTENNA__7125__CLK clknet_leaf_28_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4846__A1 _1987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5404__A _2314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4946__C _2259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3204_ _0822_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_1
XFILLER_274_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4184_ _1523_ _1688_ _1690_ _1530_ vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__o211a_1
XFILLER_267_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4962__B net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6825_ clknet_leaf_59_core_clock _0086_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[10\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5023__A1 _2301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6756_ clknet_leaf_90_core_clock _0017_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3968_ immu_0.page_table\[0\]\[1\] immu_0.page_table\[1\]\[1\] immu_0.page_table\[8\]\[1\]
+ immu_0.page_table\[9\]\[1\] _1480_ net315 vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__mux4_1
XFILLER_137_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5707_ _2709_ dmmu0.page_table\[2\]\[6\] _2702_ vssd1 vssd1 vccd1 vccd1 _2710_ sky130_fd_sc_hd__and3_1
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6687_ clknet_leaf_39_core_clock _0757_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3899_ net315 vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__clkbuf_4
XFILLER_164_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5638_ _1914_ _2217_ vssd1 vssd1 vccd1 vccd1 _2668_ sky130_fd_sc_hd__nor2_1
XFILLER_191_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5569_ _2235_ _2627_ _2630_ immu_0.page_table\[0\]\[5\] vssd1 vssd1 vccd1 vccd1 _0192_
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7308_ clknet_leaf_19_core_clock _0569_ vssd1 vssd1 vccd1 vccd1 dmmu1.long_off_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_43_core_clock clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7239_ clknet_leaf_24_core_clock _0500_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3533__S _0891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4837__A1 _1995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6129__B dmmu0.page_table\[1\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input125_A c1_o_mem_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3769__A _1334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6642__CLK clknet_leaf_56_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4591__C _2032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5984__A _1991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3576__A1 _0868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6792__CLK clknet_leaf_80_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input90_A c0_sr_bus_addr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_82_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3708__S _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5722__C1 _1911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7148__CLK clknet_leaf_34_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4828__A1 _2023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4289__C1 _1535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4766__C _2140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7298__CLK clknet_leaf_43_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6293__A3 _3058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6045__A3 _2902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5878__B _2539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5253__A1 _2233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3679__A _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4940_ _1995_ _2257_ _2260_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__a21o_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6055__A _1993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4871_ _1985_ _2195_ _2207_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__a21o_1
XFILLER_232_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3822_ _1363_ net256 vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__and2_1
X_6610_ clknet_leaf_53_core_clock _0680_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5556__A2 _2623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6541_ clknet_leaf_51_core_clock _0611_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3753_ _1326_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3618__S net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6472_ _2190_ immu_1.page_table\[8\]\[7\] _3159_ vssd1 vssd1 vccd1 vccd1 _3167_ sky130_fd_sc_hd__and3_1
X_3684_ dmmu1.page_table\[12\]\[11\] dmmu1.page_table\[13\]\[11\] _1146_ vssd1 vssd1
+ vccd1 vccd1 _1266_ sky130_fd_sc_hd__mux2_1
XFILLER_185_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5423_ net101 _2543_ vssd1 vssd1 vccd1 vccd1 _2550_ sky130_fd_sc_hd__and2_1
XFILLER_145_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3414__S1 _0863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5354_ _1929_ _2407_ vssd1 vssd1 vccd1 vccd1 _2509_ sky130_fd_sc_hd__or2_1
XFILLER_160_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6515__CLK clknet_leaf_43_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4305_ _1808_ _1809_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__xnor2_1
XFILLER_99_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5285_ _2458_ dmmu0.page_table\[14\]\[5\] _2464_ vssd1 vssd1 vccd1 vccd1 _2470_ sky130_fd_sc_hd__and3_1
XFILLER_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4819__A1 _2014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4676__C _2086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5134__A _2371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7024_ clknet_leaf_83_core_clock _0285_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4236_ immu_0.page_table\[2\]\[8\] immu_0.page_table\[3\]\[8\] _1408_ vssd1 vssd1
+ vccd1 vccd1 _1742_ sky130_fd_sc_hd__mux2_1
XFILLER_228_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6665__CLK clknet_leaf_9_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4167_ _1596_ _1674_ _1615_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__o21a_1
XFILLER_255_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_63_core_clock_A clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4098_ _1535_ _1606_ _1434_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__a21o_1
XANTENNA__5244__A1 _2211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3255__A0 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5795__A2 _2748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6808_ clknet_leaf_85_core_clock _0069_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6739_ clknet_leaf_67_core_clock _0000_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6412__B _3117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5309__A _1933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6131__C _2962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5028__B _2302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4522__A3 _1963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4586__C _2032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5044__A _1926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input242_A dcache_wb_adr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6275__A3 _3038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5483__A1 _2576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4883__A _2216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3246__A0 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6322__B _3079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5219__A _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4123__A _1462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6538__CLK clknet_leaf_48_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_core_clock core_clock vssd1 vssd1 vccd1 vccd1 clknet_0_core_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_182_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output461_A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output559_A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7434__A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5880__C _2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4513__A3 _1964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5710__A2 _2700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4269__S _1438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6688__CLK clknet_leaf_56_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5070_ _2335_ vssd1 vssd1 vccd1 vccd1 _2336_ sky130_fd_sc_hd__clkbuf_4
XFILLER_150_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5889__A _2819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4021_ _0813_ _1508_ _1515_ _1532_ vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__a31o_1
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5226__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5972_ _2799_ _2861_ vssd1 vssd1 vccd1 vccd1 _2868_ sky130_fd_sc_hd__and2_1
XFILLER_197_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4923_ _2237_ dmmu0.page_table\[0\]\[9\] _2221_ vssd1 vssd1 vccd1 vccd1 _2248_ sky130_fd_sc_hd__and3_1
XFILLER_100_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4854_ _1995_ _2195_ _2198_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__a21o_1
X_3805_ net216 _1348_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__and2_1
XFILLER_178_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4785_ _2008_ _2155_ _2160_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__a21o_1
XANTENNA__3348__S _0857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3635__S1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6524_ clknet_leaf_31_core_clock _0594_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[14\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3736_ _1302_ _1303_ _1316_ _0880_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_146_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6455_ _3156_ vssd1 vssd1 vccd1 vccd1 _3157_ sky130_fd_sc_hd__clkbuf_4
X_3667_ _1223_ _1225_ _1248_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__a21oi_1
XFILLER_173_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7344__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5790__C _2751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3399__S0 _0898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5406_ _2317_ _2439_ vssd1 vssd1 vccd1 vccd1 _2539_ sky130_fd_sc_hd__or2_4
X_6386_ _3117_ vssd1 vssd1 vccd1 vccd1 _3118_ sky130_fd_sc_hd__buf_2
XANTENNA__4504__A3 _1964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5701__A2 _2700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3598_ _0912_ _1181_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__nand2_1
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5337_ _1935_ _2497_ vssd1 vssd1 vccd1 vccd1 _2500_ sky130_fd_sc_hd__and2_1
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5268_ _2251_ _2441_ _2459_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__a21o_1
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5465__A1 _2562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5799__A _2762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4219_ net313 _1725_ vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__or2_1
X_7007_ clknet_leaf_79_core_clock _0268_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5199_ _2227_ _2409_ _2414_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__a21o_1
XFILLER_275_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3948__C_N net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5311__B _2482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5768__A2 _2729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4976__B1 _2277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5738__S _2720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6423__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5039__A _2300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input192_A c1_sr_bus_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3951__A1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3782__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6830__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input53_A c0_o_mem_long_mode vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5205__C _2411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5456__A1 _2562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6317__B _2193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5208__A1 _2240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4118__A _1442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6420__A3 _3135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7429__A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3957__A _1416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4570_ _2017_ immu_1.page_table\[14\]\[10\] _2003_ vssd1 vssd1 vccd1 vccd1 _2026_
+ sky130_fd_sc_hd__and3_1
XANTENNA__5931__A2 _2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3521_ net46 dmmu0.long_off_reg\[1\] vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__and2_1
XFILLER_155_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4788__A _2150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6240_ _2803_ _3021_ vssd1 vssd1 vccd1 vccd1 _3030_ sky130_fd_sc_hd__and2_1
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3452_ dmmu0.page_table\[0\]\[5\] dmmu0.page_table\[1\]\[5\] _0910_ vssd1 vssd1 vccd1
+ vccd1 _1040_ sky130_fd_sc_hd__mux2_1
XFILLER_226_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5695__A1 _2211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6171_ _2799_ _2983_ vssd1 vssd1 vccd1 vccd1 _2989_ sky130_fd_sc_hd__and2_1
X_3383_ dmmu0.page_table\[8\]\[2\] dmmu0.page_table\[9\]\[2\] dmmu0.page_table\[10\]\[2\]
+ dmmu0.page_table\[11\]\[2\] _0898_ _0948_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__mux4_1
XFILLER_170_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5122_ _2363_ immu_0.page_table\[13\]\[10\] _2352_ _2366_ vssd1 vssd1 vccd1 vccd1
+ _0009_ sky130_fd_sc_hd__a31o_1
XANTENNA__6239__A3 _3019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5053_ _1937_ _2322_ vssd1 vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__and2_1
XFILLER_257_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5412__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4954__C _2259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4004_ _1456_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__clkbuf_4
XFILLER_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3553__S0 _0896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6227__B _3021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6703__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6411__A3 _3115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5955_ _2856_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3867__A _1389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4906_ net100 vssd1 vssd1 vccd1 vccd1 _2235_ sky130_fd_sc_hd__buf_6
XFILLER_240_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5886_ _2777_ dmmu0.page_table\[6\]\[3\] _2814_ vssd1 vssd1 vccd1 vccd1 _2818_ sky130_fd_sc_hd__and3_1
XFILLER_178_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4837_ _1995_ _2189_ _2192_ immu_1.page_table\[1\]\[0\] vssd1 vssd1 vccd1 vccd1 _0707_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__6853__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4768_ _2134_ immu_1.page_table\[5\]\[8\] _2140_ vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__and3_1
XFILLER_217_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6507_ clknet_leaf_73_core_clock _0577_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3719_ _1207_ _1208_ _1257_ _1205_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__o211ai_1
X_4699_ _2106_ immu_1.page_table\[9\]\[2\] _2103_ vssd1 vssd1 vccd1 vccd1 _2108_ sky130_fd_sc_hd__and3_1
X_7487_ net169 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_2
XFILLER_174_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6438_ _1898_ dmmu1.page_table\[0\]\[9\] _3135_ _3147_ vssd1 vssd1 vccd1 vccd1 _0544_
+ sky130_fd_sc_hd__a31o_1
XFILLER_122_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5306__B _2367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6369_ net207 _3098_ vssd1 vssd1 vccd1 vccd1 _3107_ sky130_fd_sc_hd__and2_1
XFILLER_88_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput304 ic0_mem_data[5] vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_1
Xinput315 ic0_wb_adr[15] vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_4
Xinput326 ic0_wb_sel[0] vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_2
Xinput337 ic1_mem_data[15] vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_2
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput348 ic1_mem_data[25] vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_2
XFILLER_102_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6418__A _3136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput359 ic1_mem_data[6] vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_2
XANTENNA__5322__A _2310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6137__B dmmu0.page_table\[1\]\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5976__B _2861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6402__A3 _3116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input205_A c1_sr_bus_data_o[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3777__A _0838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5992__A _1968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3535__S0 _0865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5601__A1 _2249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4282__S _1601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5740_ immu_1.high_addr_off\[7\] _1983_ _2720_ vssd1 vssd1 vccd1 vccd1 _2728_ sky130_fd_sc_hd__mux2_1
XANTENNA__6063__A _2879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6876__CLK clknet_leaf_70_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ net710 _2687_ _1918_ _2212_ vssd1 vssd1 vccd1 vccd1 _2688_ sky130_fd_sc_hd__or4_2
XFILLER_175_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7410_ net350 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_1
X_4622_ _2019_ _2047_ _2058_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__a21o_1
XFILLER_128_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7341_ clknet_leaf_92_core_clock vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_2
XFILLER_116_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4553_ _1979_ vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__buf_6
XFILLER_156_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5407__A _1929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3504_ net152 dmmu1.long_off_reg\[2\] vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__or2_1
X_7272_ clknet_leaf_26_core_clock _0533_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_4484_ _1962_ vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__buf_2
XFILLER_143_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6223_ _1968_ _2118_ vssd1 vssd1 vccd1 vccd1 _3020_ sky130_fd_sc_hd__nor2_2
X_3435_ dmmu1.page_table\[4\]\[5\] dmmu1.page_table\[5\]\[5\] _0857_ vssd1 vssd1 vccd1
+ vccd1 _1023_ sky130_fd_sc_hd__mux2_1
XFILLER_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6154_ _2931_ vssd1 vssd1 vccd1 vccd1 _2977_ sky130_fd_sc_hd__clkbuf_4
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _0957_ _0928_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__or2_1
XFILLER_253_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _2347_ immu_0.page_table\[13\]\[2\] _2353_ _2357_ vssd1 vssd1 vccd1 vccd1
+ _0001_ sky130_fd_sc_hd__a31o_1
X_6085_ _2895_ _2923_ vssd1 vssd1 vccd1 vccd1 _2937_ sky130_fd_sc_hd__and2_1
XFILLER_253_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6238__A _2801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ _0875_ _0880_ _0889_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__and3_2
XANTENNA__4684__C _2086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5142__A _2371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ net93 vssd1 vssd1 vccd1 vccd1 _2314_ sky130_fd_sc_hd__buf_4
XFILLER_38_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6987_ clknet_leaf_7_core_clock _0248_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3603__B1 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5938_ net95 _2829_ _2847_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__a21o_1
XFILLER_278_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5869_ _2805_ dmmu1.page_table\[15\]\[9\] _2787_ _2807_ vssd1 vssd1 vccd1 vccd1 _0315_
+ sky130_fd_sc_hd__a31o_1
XFILLER_278_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5371__A3 _2510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5317__A _1942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4859__C _2197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5659__A1 _2245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7181__CLK clknet_leaf_29_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input155_A c1_o_mem_high_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput101 c0_sr_bus_data_o[6] vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__buf_4
XFILLER_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput112 c1_o_instr_long_addr[2] vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_2
Xinput123 c1_o_mem_addr[14] vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_4
XFILLER_48_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput134 c1_o_mem_data[0] vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_2
Xinput145 c1_o_mem_data[5] vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_2
XFILLER_130_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6148__A _2971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6084__A1 _2932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput156 c1_o_mem_high_addr[6] vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput167 c1_o_req_addr[12] vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input322_A ic0_wb_adr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput178 c1_o_req_addr[8] vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput189 c1_sr_bus_addr[2] vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_4
XFILLER_236_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5831__A1 _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input16_A c0_o_mem_addr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4891__A _2223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6899__CLK clknet_leaf_76_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5898__A1 _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3954__B _1416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6330__B _3079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5362__A3 _2510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput608 net608 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[0] sky130_fd_sc_hd__buf_2
XFILLER_125_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput619 net619 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[5] sky130_fd_sc_hd__buf_2
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output541_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output639_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7442__A net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3970__A _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4322__A1 _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3220_ net215 _0824_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__and2_1
XFILLER_97_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4873__A2 _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6058__A _2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5897__A _2819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5822__A1 _2239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6910_ clknet_leaf_76_core_clock _0171_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_282_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6841_ clknet_leaf_68_core_clock _0102_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_68_core_clock_A clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4389__A1 _1890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6772_ clknet_leaf_91_core_clock _0033_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[9\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3210__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3984_ _1487_ _1492_ _1495_ _1496_ _0812_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__o221a_1
XFILLER_250_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5723_ net191 vssd1 vssd1 vccd1 vccd1 _2718_ sky130_fd_sc_hd__inv_2
XFILLER_188_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5654_ _2666_ dmmu0.page_table\[11\]\[6\] _2671_ vssd1 vssd1 vccd1 vccd1 _2678_ sky130_fd_sc_hd__and3_1
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4605_ _2048_ vssd1 vssd1 vccd1 vccd1 _2049_ sky130_fd_sc_hd__buf_2
XFILLER_148_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6240__B _3021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5585_ _2473_ dmmu0.page_table\[12\]\[3\] _2634_ vssd1 vssd1 vccd1 vccd1 _2638_ sky130_fd_sc_hd__and3_1
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4010__B1 _1521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4536_ _2001_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__clkbuf_4
XFILLER_190_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_core_clock clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7255_ clknet_leaf_21_core_clock _0516_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5105__A3 _2353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4467_ net104 vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__buf_6
XANTENNA__3880__A _1398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4313__A1 _1523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6206_ _2994_ dmmu1.page_table\[7\]\[6\] _3000_ _3009_ vssd1 vssd1 vccd1 vccd1 _0450_
+ sky130_fd_sc_hd__a31o_1
XFILLER_89_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3418_ _0995_ net124 vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__and2b_2
X_4398_ _1896_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__buf_6
X_7186_ clknet_leaf_16_core_clock _0447_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4864__A2 _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input8_A c0_o_instr_long_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3349_ _0863_ _0940_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__or2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6137_ _2845_ dmmu0.page_table\[1\]\[5\] _2962_ vssd1 vssd1 vccd1 vccd1 _2968_ sky130_fd_sc_hd__and3_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6066__A1 _2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6068_ _2914_ dmmu1.page_table\[10\]\[2\] _2922_ _2927_ vssd1 vssd1 vccd1 vccd1 _0394_
+ sky130_fd_sc_hd__a31o_1
XFILLER_277_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4616__A2 _2047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5019_ _2301_ immu_0.page_table\[15\]\[2\] _2298_ _2304_ vssd1 vssd1 vccd1 vccd1
+ _0777_ sky130_fd_sc_hd__a31o_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5600__A _2640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_72_core_clock clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6431__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4001__B1 _1512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4589__C _2032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5047__A _1928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4552__A1 _2012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_70_core_clock_A clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_5_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input272_A dcache_wb_sel[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6571__CLK clknet_leaf_46_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4886__A _2212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3790__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4304__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5213__C _2411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4607__A2 _2047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5804__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5280__A2 _2462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7437__A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3965__A _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6341__A _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4791__A1 _2014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6914__CLK clknet_leaf_79_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4543__A1 _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput405 net405 vssd1 vssd1 vccd1 vccd1 c0_clk sky130_fd_sc_hd__clkbuf_1
X_5370_ _1942_ _2512_ vssd1 vssd1 vccd1 vccd1 _2519_ sky130_fd_sc_hd__and2_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput416 net416 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[13] sky130_fd_sc_hd__buf_2
Xoutput427 net427 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[9] sky130_fd_sc_hd__buf_2
XFILLER_126_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4321_ _1581_ _1825_ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__or2_1
XFILLER_113_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput438 net438 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[18] sky130_fd_sc_hd__buf_2
XANTENNA__6487__S _3172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4796__A _2105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4387__A2_N _1889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput449 net449 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[28] sky130_fd_sc_hd__buf_2
XFILLER_4_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3729__S0 _1146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7040_ clknet_leaf_12_core_clock _0301_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_4252_ net114 immu_1.high_addr_off\[4\] vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__or2_1
XANTENNA__4846__A2 _2189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3203_ net222 _0819_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__and2_1
XANTENNA__5404__B _2527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4183_ _1442_ _1689_ vssd1 vssd1 vccd1 vccd1 _1690_ sky130_fd_sc_hd__or2_1
XFILLER_255_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3205__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4962__C net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3901__S0 _1407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3282__A1 _0855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6824_ clknet_leaf_59_core_clock _0085_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[10\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6755_ clknet_leaf_89_core_clock _0016_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3967_ _1472_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__buf_6
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5706_ _2681_ vssd1 vssd1 vccd1 vccd1 _2709_ sky130_fd_sc_hd__clkbuf_4
XFILLER_259_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6686_ clknet_leaf_56_core_clock _0756_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3898_ _1409_ _1411_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__or2_1
XANTENNA__6594__CLK clknet_leaf_54_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5637_ _2253_ _2649_ _2667_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__a21o_1
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3968__S0 _1480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5568_ _2232_ _2627_ _2630_ immu_0.page_table\[0\]\[4\] vssd1 vssd1 vccd1 vccd1 _0191_
+ sky130_fd_sc_hd__o22a_1
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7307_ clknet_leaf_19_core_clock _0568_ vssd1 vssd1 vccd1 vccd1 dmmu1.long_off_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4519_ _1976_ dmmu1.page_table\[14\]\[9\] _1964_ _1988_ vssd1 vssd1 vccd1 vccd1 _0593_
+ sky130_fd_sc_hd__a31o_1
XFILLER_144_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5499_ net98 _2593_ vssd1 vssd1 vccd1 vccd1 _2596_ sky130_fd_sc_hd__and2_1
XFILLER_78_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7238_ clknet_leaf_20_core_clock _0499_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4837__A2 _2189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7169_ clknet_leaf_3_core_clock _0430_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6039__A1 _2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6129__C _2962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4872__C _2197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5330__A _1926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input118_A c1_o_mem_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6211__A1 _3010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6937__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6161__A _2879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input83_A c0_sr_bus_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4525__A1 _1976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3733__C1 _0854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3724__S _1146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5505__A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4828__A2 _2172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4782__C _2157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5240__A _2215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5253__A2 _2442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4870_ _2204_ immu_1.page_table\[3\]\[8\] _2197_ vssd1 vssd1 vccd1 vccd1 _2207_ sky130_fd_sc_hd__and3_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6202__A1 _2994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3821_ inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__buf_4
XFILLER_60_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4290__S _1425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6071__A _2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6540_ clknet_leaf_51_core_clock _0610_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3752_ net146 net41 _1322_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__mux2_2
XFILLER_146_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6471_ _1981_ _3157_ _3166_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__a21o_1
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3683_ _0869_ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__nor2_1
XANTENNA__5308__A3 _2480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4516__A1 _1976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5422_ _2546_ immu_0.page_table\[6\]\[5\] _2541_ _2549_ vssd1 vssd1 vccd1 vccd1 _0126_
+ sky130_fd_sc_hd__a31o_1
XFILLER_133_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5353_ _2503_ immu_0.page_table\[9\]\[10\] _2494_ _2508_ vssd1 vssd1 vccd1 vccd1
+ _0098_ sky130_fd_sc_hd__a31o_1
XANTENNA__6269__A1 _3042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4304_ net114 immu_1.high_addr_off\[4\] _1759_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__a21o_1
X_5284_ _2233_ _2462_ _2469_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__a21o_1
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4819__A2 _2172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7023_ clknet_leaf_82_core_clock _0284_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4235_ immu_0.page_table\[0\]\[8\] immu_0.page_table\[1\]\[8\] _1409_ vssd1 vssd1
+ vccd1 vccd1 _1741_ sky130_fd_sc_hd__mux2_1
XFILLER_247_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4166_ net111 immu_1.high_addr_off\[1\] vssd1 vssd1 vccd1 vccd1 _1674_ sky130_fd_sc_hd__nor2_1
XFILLER_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6246__A _2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5788__C _2751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4097_ immu_0.page_table\[8\]\[5\] immu_0.page_table\[9\]\[5\] immu_0.page_table\[10\]\[5\]
+ immu_0.page_table\[11\]\[5\] _1601_ _1420_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__mux4_1
XANTENNA__5150__A _2370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5244__A2 _2442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6807_ clknet_leaf_82_core_clock _0068_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4999_ _2284_ immu_1.page_table\[15\]\[7\] _2282_ vssd1 vssd1 vccd1 vccd1 _2291_
+ sky130_fd_sc_hd__and3_1
XFILLER_196_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4755__A1 _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6738_ clknet_leaf_66_core_clock _0808_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5309__B _2482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6669_ clknet_leaf_3_core_clock _0739_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4507__A1 _1976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3715__C1 _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5180__A1 _2245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input235_A dcache_wb_adr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6156__A _2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5698__C _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6432__A1 _1898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input402_A inner_wb_i_dat[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4994__A1 _1977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7115__CLK clknet_leaf_30_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4746__A1 _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4123__B _1625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5171__A1 _2233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output454_A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3454__S _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7450__A net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4020_ _1516_ _1522_ _1528_ _1531_ _0812_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__o221a_1
XFILLER_284_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5226__A2 _2430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5971_ _2561_ vssd1 vssd1 vccd1 vccd1 _2867_ sky130_fd_sc_hd__buf_4
XFILLER_213_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4985__A1 _1995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4922_ _1948_ vssd1 vssd1 vccd1 vccd1 _2247_ sky130_fd_sc_hd__buf_4
XFILLER_240_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4853_ _2182_ immu_1.page_table\[3\]\[0\] _2197_ vssd1 vssd1 vccd1 vccd1 _2198_ sky130_fd_sc_hd__and3_1
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5529__A3 _2607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3629__S _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3804_ _1353_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4737__A1 _2016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4784_ _2150_ immu_1.page_table\[4\]\[2\] _2157_ vssd1 vssd1 vccd1 vccd1 _2160_ sky130_fd_sc_hd__and3_1
XFILLER_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6523_ clknet_leaf_44_core_clock _0593_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[14\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3735_ _1307_ _1309_ _1315_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__a21oi_4
XFILLER_118_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6454_ _1999_ _2978_ vssd1 vssd1 vccd1 vccd1 _3156_ sky130_fd_sc_hd__nor2_1
XFILLER_146_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3666_ _1222_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__inv_2
XFILLER_134_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5405_ _2531_ immu_0.page_table\[7\]\[10\] _2524_ _2538_ vssd1 vssd1 vccd1 vccd1
+ _0120_ sky130_fd_sc_hd__a31o_1
XANTENNA__3399__S1 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6385_ _2784_ _2187_ vssd1 vssd1 vccd1 vccd1 _3117_ sky130_fd_sc_hd__nor2_1
XANTENNA__6632__CLK clknet_leaf_41_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3597_ dmmu0.page_table\[6\]\[9\] dmmu0.page_table\[7\]\[9\] _1169_ vssd1 vssd1 vccd1
+ vccd1 _1181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5336_ _2489_ immu_0.page_table\[9\]\[2\] _2495_ _2499_ vssd1 vssd1 vccd1 vccd1 _0090_
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4984__A _2262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5267_ _2458_ dmmu0.page_table\[7\]\[11\] _2444_ vssd1 vssd1 vccd1 vccd1 _2459_ sky130_fd_sc_hd__and3_1
XFILLER_102_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7006_ clknet_leaf_80_core_clock _0267_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4122__C1 _1553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4218_ immu_0.page_table\[8\]\[7\] immu_0.page_table\[9\]\[7\] net312 vssd1 vssd1
+ vccd1 vccd1 _1725_ sky130_fd_sc_hd__mux2_1
X_5198_ _2400_ dmmu0.page_table\[8\]\[2\] _2411_ vssd1 vssd1 vccd1 vccd1 _2414_ sky130_fd_sc_hd__and3_1
XFILLER_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4149_ _1447_ _1656_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__or2_1
XFILLER_228_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7138__CLK clknet_leaf_28_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4976__A1 _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6423__B _3137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4224__A inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input185_A c1_sr_bus_addr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3782__B _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4597__C _2032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5055__A _1940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input352_A ic1_mem_data[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input46_A c0_o_mem_high_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4894__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3303__A _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5208__A2 _2409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4967__B2 immu_1.page_table\[0\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6505__CLK clknet_leaf_62_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6333__B _3079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3449__S _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3973__A _1447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6655__CLK clknet_leaf_39_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7445__A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3520_ net47 dmmu0.long_off_reg\[2\] vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__nor2_1
XANTENNA__5891__C _2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3451_ _0909_ _1036_ _1038_ _0906_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__o211a_1
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5695__A2 _2700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6170_ _2977_ dmmu1.page_table\[8\]\[4\] _2981_ _2988_ vssd1 vssd1 vccd1 vccd1 _0435_
+ sky130_fd_sc_hd__a31o_1
X_3382_ dmmu0.page_table\[0\]\[2\] dmmu0.page_table\[1\]\[2\] dmmu0.page_table\[2\]\[2\]
+ dmmu0.page_table\[3\]\[2\] _0898_ _0948_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__mux4_1
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5121_ _2314_ _2355_ vssd1 vssd1 vccd1 vccd1 _2366_ sky130_fd_sc_hd__and2_1
XFILLER_97_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6495__S _3172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3912__S _1425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5052_ _2316_ immu_0.page_table\[14\]\[3\] _2320_ _2325_ vssd1 vssd1 vccd1 vccd1
+ _0789_ sky130_fd_sc_hd__a31o_1
XFILLER_111_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5412__B _2543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4003_ _1434_ _1509_ _1513_ _1514_ vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__a211o_1
XFILLER_284_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3553__S1 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5954_ dmmu0.long_off_reg\[7\] _1944_ _2848_ vssd1 vssd1 vccd1 vccd1 _2856_ sky130_fd_sc_hd__mux2_1
XFILLER_225_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4905_ _2233_ _2219_ _2234_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__a21o_1
XFILLER_178_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5885_ _2226_ _2812_ _2817_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__a21o_1
XANTENNA__3359__S _0900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4836_ _2191_ vssd1 vssd1 vccd1 vccd1 _2192_ sky130_fd_sc_hd__clkbuf_4
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_0_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_193_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5383__A1 _2517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4767_ _2019_ _2138_ _2148_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__a21o_1
XANTENNA__3883__A _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6506_ clknet_leaf_68_core_clock _0576_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3394__B1 _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3718_ _0957_ _1283_ _1284_ _1298_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__a31o_1
X_7486_ net168 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__buf_2
X_4698_ _2006_ _2101_ _2107_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__a21o_1
XFILLER_112_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5135__A1 _2227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6437_ net209 _3137_ vssd1 vssd1 vccd1 vccd1 _3147_ sky130_fd_sc_hd__and2_1
XFILLER_146_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3649_ dmmu0.page_table\[0\]\[11\] dmmu0.page_table\[1\]\[11\] _0895_ vssd1 vssd1
+ vccd1 vccd1 _1231_ sky130_fd_sc_hd__mux2_1
XFILLER_283_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_75_core_clock_A clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_136_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6368_ _3101_ dmmu1.page_table\[2\]\[6\] _3096_ _3106_ vssd1 vssd1 vccd1 vccd1 _0515_
+ sky130_fd_sc_hd__a31o_1
XFILLER_121_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5319_ _2300_ vssd1 vssd1 vccd1 vccd1 _2489_ sky130_fd_sc_hd__buf_4
XFILLER_276_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6299_ _3053_ dmmu1.page_table\[4\]\[4\] _3058_ _3065_ vssd1 vssd1 vccd1 vccd1 _0487_
+ sky130_fd_sc_hd__a31o_1
Xinput305 ic0_mem_data[6] vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_1
Xinput316 ic0_wb_adr[1] vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_2
XFILLER_29_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput327 ic0_wb_sel[1] vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_2
XFILLER_48_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput338 ic1_mem_data[16] vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__buf_2
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput349 ic1_mem_data[26] vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_2
XFILLER_248_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5322__B _2482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4219__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6137__C _2962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6528__CLK clknet_leaf_41_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4949__A1 _1977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input100_A c0_sr_bus_data_o[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3777__B _1168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3621__A1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6166__A3 _2981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5992__B _2045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3385__B1 _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5513__A _2561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6328__B _3079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3535__S1 _0863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5886__C _2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4790__C _2157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6063__B _2924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ net86 vssd1 vssd1 vccd1 vccd1 _2687_ sky130_fd_sc_hd__clkinv_2
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4621_ _2054_ immu_1.page_table\[12\]\[7\] _2049_ vssd1 vssd1 vccd1 vccd1 _2058_
+ sky130_fd_sc_hd__and3_1
XFILLER_175_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4799__A _2166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3907__S _1408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3376__B1 _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4552_ _2012_ _2002_ _2013_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__a21o_1
XFILLER_237_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3471__S0 _0858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_core_clock clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5407__B _2539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3503_ net152 dmmu1.long_off_reg\[2\] vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__nand2_1
X_7271_ clknet_leaf_25_core_clock _0532_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4483_ _1958_ _1961_ vssd1 vssd1 vccd1 vccd1 _1962_ sky130_fd_sc_hd__or2_1
XFILLER_171_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3208__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6222_ _3018_ vssd1 vssd1 vccd1 vccd1 _3019_ sky130_fd_sc_hd__buf_4
X_3434_ dmmu1.page_table\[6\]\[5\] dmmu1.page_table\[7\]\[5\] _0865_ vssd1 vssd1 vccd1
+ vccd1 _1022_ sky130_fd_sc_hd__mux2_1
XFILLER_171_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ net95 _2959_ _2976_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__a21o_1
XFILLER_258_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _0927_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__clkbuf_4
XFILLER_106_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5423__A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _1933_ _2355_ vssd1 vssd1 vccd1 vccd1 _2357_ sky130_fd_sc_hd__and2_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _2932_ dmmu1.page_table\[10\]\[9\] _2922_ _2936_ vssd1 vssd1 vccd1 vccd1 _0401_
+ sky130_fd_sc_hd__a31o_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6238__B _3021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _0881_ _0883_ _0885_ _0888_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__a31o_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5035_ _2301_ immu_0.page_table\[15\]\[9\] _2298_ _2313_ vssd1 vssd1 vccd1 vccd1
+ _0784_ sky130_fd_sc_hd__a31o_1
XFILLER_272_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5796__C _2751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6820__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6986_ clknet_leaf_7_core_clock _0247_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_280_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6396__A3 _3116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5937_ _2845_ dmmu0.page_table\[5\]\[12\] _2831_ vssd1 vssd1 vccd1 vccd1 _2847_ sky130_fd_sc_hd__and3_1
XANTENNA__3603__A1 _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_62_core_clock clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5868_ _1987_ _2789_ vssd1 vssd1 vccd1 vccd1 _2807_ sky130_fd_sc_hd__and2_1
XFILLER_221_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4819_ _2014_ _2172_ _2180_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__a21o_1
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5799_ _2762_ dmmu0.page_table\[13\]\[10\] _2750_ vssd1 vssd1 vccd1 vccd1 _2763_
+ sky130_fd_sc_hd__and3_1
XANTENNA__3367__B1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4502__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5317__B _2482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3382__A3 dmmu0.page_table\[3\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7469_ net393 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5659__A2 _2669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3552__S _0918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5333__A _1928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput102 c0_sr_bus_data_o[7] vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__buf_4
XFILLER_248_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput113 c1_o_instr_long_addr[3] vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_2
Xinput124 c1_o_mem_addr[15] vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput135 c1_o_mem_data[10] vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input148_A c1_o_mem_data[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput146 c1_o_mem_data[6] vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_2
Xinput157 c1_o_mem_high_addr[7] vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput168 c1_o_req_addr[13] vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput179 c1_o_req_addr[9] vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4095__A1 _1479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input315_A ic0_wb_adr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3788__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5595__A1 _2243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5347__A1 _2503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5898__A2 _2812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4412__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput609 net609 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[10] sky130_fd_sc_hd__buf_2
XFILLER_165_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5942__S _2848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6339__A _2891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3462__S _0900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5243__A _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6058__B _2081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_255_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6843__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_1_0_0_core_clock_A clknet_0_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6840_ clknet_leaf_69_core_clock _0101_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6771_ clknet_leaf_89_core_clock _0032_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[9\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5586__A1 _2230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6993__CLK clknet_leaf_5_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3983_ _1442_ vssd1 vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__buf_4
XFILLER_250_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3210__B _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0_core_clock clknet_1_1_1_core_clock vssd1 vssd1 vccd1 vccd1 clknet_2_3_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__5050__A3 _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5722_ _1579_ net379 _2717_ _1911_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__o211a_1
XFILLER_148_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5338__A1 _2489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5653_ _2236_ _2669_ _2677_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__a21o_1
XFILLER_148_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4604_ _1999_ _2045_ vssd1 vssd1 vccd1 vccd1 _2048_ sky130_fd_sc_hd__or2_1
XFILLER_191_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5584_ _2227_ _2632_ _2637_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__a21o_1
XANTENNA__4010__A1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4535_ _1961_ _2000_ vssd1 vssd1 vccd1 vccd1 _2001_ sky130_fd_sc_hd__nor2_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7254_ clknet_leaf_21_core_clock _0515_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4466_ _1939_ immu_0.page_table\[11\]\[8\] _1924_ _1947_ vssd1 vssd1 vccd1 vccd1
+ _0581_ sky130_fd_sc_hd__a31o_1
XFILLER_131_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6205_ _2801_ _3002_ vssd1 vssd1 vccd1 vccd1 _3009_ sky130_fd_sc_hd__and2_1
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5510__A1 _2588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3417_ _0995_ _0996_ _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__o21a_2
X_7185_ clknet_leaf_13_core_clock _0446_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4397_ net710 vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__inv_2
XANTENNA__5153__A _2384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _2232_ _2960_ _2967_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__a21o_1
X_3348_ dmmu1.page_table\[4\]\[1\] dmmu1.page_table\[5\]\[1\] _0857_ vssd1 vssd1 vccd1
+ vccd1 _0940_ sky130_fd_sc_hd__mux2_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6067_ _2793_ _2924_ vssd1 vssd1 vccd1 vccd1 _2927_ sky130_fd_sc_hd__and2_1
XFILLER_280_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3279_ _0871_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__buf_4
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4077__A1 _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5018_ _1933_ _2302_ vssd1 vssd1 vccd1 vccd1 _2304_ sky130_fd_sc_hd__and2_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6969_ clknet_leaf_86_core_clock _0230_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6431__B _3137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5328__A _1929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4001__A1 _1424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5047__B _2322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6716__CLK clknet_leaf_62_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4552__A2 _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3760__A0 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input265_A dcache_wb_o_dat[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4886__B _2215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3790__B _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6159__A _1968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6866__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5063__A _2312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5998__A _2561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5804__A2 _2747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5568__A1 _2232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5032__A3 _2298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6341__B _3079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4791__A2 _2155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3457__S _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5238__A _2217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4142__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3426__S0 _0897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4543__A2 _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5740__A1 _1983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput406 net406 vssd1 vssd1 vccd1 vccd1 c0_disable sky130_fd_sc_hd__buf_2
XANTENNA__7453__A net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput417 net417 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[14] sky130_fd_sc_hd__buf_2
X_4320_ immu_1.page_table\[0\]\[9\] immu_1.page_table\[1\]\[9\] _1493_ vssd1 vssd1
+ vccd1 vccd1 _1825_ sky130_fd_sc_hd__mux2_1
Xoutput428 net428 vssd1 vssd1 vccd1 vccd1 c0_i_mem_exception sky130_fd_sc_hd__buf_2
XFILLER_141_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput439 net439 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[19] sky130_fd_sc_hd__buf_2
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4251_ _1676_ _1682_ _1683_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__o21ai_1
XANTENNA__3729__S1 _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6069__A _2795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3202_ _0821_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_1
XFILLER_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4182_ immu_1.page_table\[0\]\[7\] immu_1.page_table\[1\]\[7\] _1443_ vssd1 vssd1
+ vccd1 vccd1 _1689_ sky130_fd_sc_hd__mux2_1
XFILLER_67_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3205__B _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7021__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4962__D net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3901__S1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3221__A _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6823_ clknet_leaf_74_core_clock _0084_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7171__CLK clknet_leaf_33_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5023__A3 _2298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6754_ clknet_leaf_89_core_clock _0015_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3966_ _1432_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5705_ _2236_ _2700_ _2708_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__a21o_1
XFILLER_148_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6685_ clknet_leaf_57_core_clock _0755_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3897_ _1410_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5148__A _2371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5636_ _2666_ dmmu0.page_table\[15\]\[12\] _2651_ vssd1 vssd1 vccd1 vccd1 _2667_
+ sky130_fd_sc_hd__and3_1
XANTENNA__3990__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_14_core_clock_A clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4987__A _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5567_ _2229_ _2627_ _2630_ immu_0.page_table\[0\]\[3\] vssd1 vssd1 vccd1 vccd1 _0190_
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3968__S1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7306_ clknet_leaf_18_core_clock _0567_ vssd1 vssd1 vccd1 vccd1 dmmu1.long_off_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4518_ _1987_ _1970_ vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__and2_1
X_5498_ _2588_ immu_0.page_table\[3\]\[2\] _2591_ _2595_ vssd1 vssd1 vccd1 vccd1 _0156_
+ sky130_fd_sc_hd__a31o_1
XFILLER_132_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7237_ clknet_leaf_21_core_clock _0498_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4449_ _1935_ _1931_ vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__and2_1
XANTENNA__4298__A1 _1535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7168_ clknet_leaf_4_core_clock _0429_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6119_ _1991_ _2943_ vssd1 vssd1 vccd1 vccd1 _2957_ sky130_fd_sc_hd__and2_1
XFILLER_258_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7099_ clknet_leaf_32_core_clock _0360_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4227__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5970__A1 _2805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6161__B _2983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3277__S _0858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input382_A ic1_wb_stb vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3408__S0 _0891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input76_A c0_sr_bus_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5722__A1 _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5505__B _2593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4289__A1 _1570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3306__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7044__CLK clknet_leaf_4_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5521__A _1922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5789__A1 _2235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7194__CLK clknet_leaf_27_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7448__A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3976__A _1451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3820_ _1362_ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__clkbuf_1
XFILLER_260_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_3_0_core_clock_A clknet_2_1_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_260_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6352__A _2784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3751_ _1325_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_1
XANTENNA__6071__B _2924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6470_ _2190_ immu_1.page_table\[8\]\[6\] _3159_ vssd1 vssd1 vccd1 vccd1 _3166_ sky130_fd_sc_hd__and3_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3682_ dmmu1.page_table\[14\]\[11\] dmmu1.page_table\[15\]\[11\] _1146_ vssd1 vssd1
+ vccd1 vccd1 _1264_ sky130_fd_sc_hd__mux2_1
XFILLER_118_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_5_core_clock_A clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5421_ net100 _2543_ vssd1 vssd1 vccd1 vccd1 _2549_ sky130_fd_sc_hd__and2_1
XANTENNA__4072__S0 _1439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5352_ _2314_ _2497_ vssd1 vssd1 vccd1 vccd1 _2508_ sky130_fd_sc_hd__and2_1
XFILLER_99_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4303_ _1806_ _1807_ vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__or2b_1
X_5283_ _2458_ dmmu0.page_table\[14\]\[4\] _2464_ vssd1 vssd1 vccd1 vccd1 _2469_ sky130_fd_sc_hd__and3_1
XFILLER_245_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3216__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7022_ clknet_leaf_83_core_clock _0283_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5134__C _2373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4234_ _1570_ _1737_ _1739_ _1479_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__o211a_1
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4165_ _1441_ _1663_ _1672_ vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__and3_1
XANTENNA__5431__A _2314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6246__B _3020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4096_ immu_0.page_table\[12\]\[5\] immu_0.page_table\[13\]\[5\] immu_0.page_table\[14\]\[5\]
+ immu_0.page_table\[15\]\[5\] _1409_ _1570_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__mux4_1
XFILLER_255_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6561__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3660__C1 _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3886__A _1402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6806_ clknet_leaf_84_core_clock _0067_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6262__A _2793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4998_ _1981_ _2280_ _2290_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__a21o_1
XFILLER_211_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6737_ clknet_leaf_66_core_clock _0807_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[12\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5952__A1 _1942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4755__A2 _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3949_ net369 _1461_ _1462_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__a21o_1
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6668_ clknet_leaf_5_core_clock _0738_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5619_ _2655_ dmmu0.page_table\[15\]\[4\] _2652_ vssd1 vssd1 vccd1 vccd1 _2658_ sky130_fd_sc_hd__and3_1
X_6599_ clknet_leaf_56_core_clock _0669_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4063__S0 _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5606__A _2217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5180__A2 _2390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7067__CLK clknet_leaf_5_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5483__A3 _2574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3560__S _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6437__A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5341__A _1940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input130_A c1_o_mem_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input228_A dcache_mem_o_data[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6904__CLK clknet_leaf_79_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4994__A2 _2280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_82_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__C1 _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4391__S _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6196__A1 _2994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4404__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4420__A _1897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5171__A2 _2390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5950__S _2848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output447_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6120__A1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6347__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5889__C _2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5970_ _2805_ dmmu1.page_table\[13\]\[4\] _2859_ _2866_ vssd1 vssd1 vccd1 vccd1 _0357_
+ sky130_fd_sc_hd__a31o_1
XFILLER_18_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4921_ _2245_ _2219_ _2246_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__a21o_1
XFILLER_280_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4985__A2 _2280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6187__A1 _2994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4852_ _2196_ vssd1 vssd1 vccd1 vccd1 _2197_ sky130_fd_sc_hd__buf_2
XFILLER_205_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3803_ net215 _1348_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__and2_1
XANTENNA__4198__B1 _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4737__A2 _2120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4783_ _2006_ _2155_ _2159_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__a21o_1
XFILLER_193_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6522_ clknet_leaf_43_core_clock _0592_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[14\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3734_ _0872_ _1310_ _1314_ _0874_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__a211oi_2
XFILLER_220_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6453_ net710 _3155_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__nor2_1
X_3665_ _0921_ _1242_ _1246_ _0929_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__o31a_1
XFILLER_118_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5404_ _2314_ _2527_ vssd1 vssd1 vccd1 vccd1 _2538_ sky130_fd_sc_hd__and2_1
XFILLER_256_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6384_ _3115_ vssd1 vssd1 vccd1 vccd1 _3116_ sky130_fd_sc_hd__clkbuf_4
X_3596_ _0908_ _1179_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__nand2_1
X_5335_ _1933_ _2497_ vssd1 vssd1 vccd1 vccd1 _2499_ sky130_fd_sc_hd__and2_1
XFILLER_114_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5266_ _2370_ vssd1 vssd1 vccd1 vccd1 _2458_ sky130_fd_sc_hd__clkbuf_4
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7005_ clknet_leaf_36_core_clock _0266_ vssd1 vssd1 vccd1 vccd1 immu_1.high_addr_off\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_275_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5465__A3 _2574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4217_ immu_0.page_table\[10\]\[7\] immu_0.page_table\[11\]\[7\] _1407_ vssd1 vssd1
+ vccd1 vccd1 _1724_ sky130_fd_sc_hd__mux2_1
XFILLER_102_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5799__C _2750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6257__A _2879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5197_ _2224_ _2409_ _2413_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__a21o_1
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4673__A1 _2010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4148_ immu_1.page_table\[14\]\[6\] immu_1.page_table\[15\]\[6\] _1437_ vssd1 vssd1
+ vccd1 vccd1 _1656_ sky130_fd_sc_hd__mux2_1
XFILLER_228_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4079_ immu_1.page_table\[4\]\[4\] immu_1.page_table\[5\]\[4\] _1524_ vssd1 vssd1
+ vccd1 vccd1 _1589_ sky130_fd_sc_hd__mux2_1
XFILLER_243_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4976__A2 _2274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6178__A1 _2977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5925__A1 _2239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4224__B _1706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3951__A3 _1436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3555__S _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input178_A c1_o_req_addr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5055__B _2322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input345_A ic1_mem_data[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5456__A3 _2557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_A c0_o_mem_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6167__A _2795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5071__A _1926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7232__CLK clknet_leaf_27_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3973__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_core_clock clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5246__A _2447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4788__C _2157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3450_ _0948_ _1037_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__or2_1
XFILLER_128_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3381_ _0958_ _0969_ _0971_ _0906_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__o31a_1
XFILLER_226_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5680__S _2690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7461__A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5120_ _2363_ immu_0.page_table\[13\]\[9\] _2353_ _2365_ vssd1 vssd1 vccd1 vccd1
+ _0008_ sky130_fd_sc_hd__a31o_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4104__B1 _1360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5051_ _1935_ _2322_ vssd1 vssd1 vccd1 vccd1 _2325_ sky130_fd_sc_hd__and2_1
XFILLER_284_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6077__A _2801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4002_ _1432_ _1410_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__nand2_1
XFILLER_272_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5953_ _2855_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_280_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4904_ _2204_ dmmu0.page_table\[0\]\[4\] _2221_ vssd1 vssd1 vccd1 vccd1 _2234_ sky130_fd_sc_hd__and3_1
XANTENNA__4325__A _1363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5884_ _2777_ dmmu0.page_table\[6\]\[2\] _2814_ vssd1 vssd1 vccd1 vccd1 _2817_ sky130_fd_sc_hd__and3_1
XFILLER_240_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4835_ _2190_ _2188_ vssd1 vssd1 vccd1 vccd1 _2191_ sky130_fd_sc_hd__nand2_1
XFILLER_178_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4766_ _2134_ immu_1.page_table\[5\]\[7\] _2140_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__and3_1
XFILLER_119_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3394__A1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3717_ _1291_ _1297_ _0929_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__and3b_1
X_6505_ clknet_leaf_62_core_clock _0575_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_267_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7485_ net167 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__buf_2
X_4697_ _2106_ immu_1.page_table\[9\]\[1\] _2103_ vssd1 vssd1 vccd1 vccd1 _2107_ sky130_fd_sc_hd__and3_1
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3375__S _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4060__A _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6436_ _1898_ dmmu1.page_table\[0\]\[8\] _3135_ _3146_ vssd1 vssd1 vccd1 vccd1 _0543_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__5135__A2 _2369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3648_ dmmu0.page_table\[2\]\[11\] dmmu0.page_table\[3\]\[11\] _1169_ vssd1 vssd1
+ vccd1 vccd1 _1230_ sky130_fd_sc_hd__mux2_1
XFILLER_161_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4995__A _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6367_ net206 _3098_ vssd1 vssd1 vccd1 vccd1 _3106_ sky130_fd_sc_hd__and2_1
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3579_ net154 dmmu1.long_off_reg\[4\] vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__nand2_1
XFILLER_283_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5318_ _2363_ immu_0.page_table\[10\]\[6\] _2480_ _2488_ vssd1 vssd1 vccd1 vccd1
+ _0083_ sky130_fd_sc_hd__a31o_1
X_6298_ net204 _3060_ vssd1 vssd1 vccd1 vccd1 _3065_ sky130_fd_sc_hd__and2_1
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput306 ic0_mem_data[7] vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput317 ic0_wb_adr[2] vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_2
Xinput328 ic0_wb_stb vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_2
X_5249_ _2227_ _2442_ _2449_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__a21o_1
Xinput339 ic1_mem_data[17] vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_2
XANTENNA__7105__CLK clknet_leaf_35_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4646__A1 _2012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3404__A _0839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_91_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4949__A2 _2257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3777__C _1211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6450__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input295_A ic0_mem_data[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3385__A1 _0918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5066__A _2314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6323__A1 _3069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4637__A1 _1996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5062__A1 _2316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6622__CLK clknet_leaf_62_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7456__A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4620_ _2016_ _2047_ _2057_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__a21o_1
XANTENNA__3376__A1 _0881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4551_ _1910_ immu_1.page_table\[14\]\[4\] _2004_ vssd1 vssd1 vccd1 vccd1 _2013_
+ sky130_fd_sc_hd__and3_1
XFILLER_128_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3471__S1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3502_ net106 net158 _0835_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__o21a_2
X_7270_ clknet_leaf_25_core_clock _0531_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6314__A1 _3069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4482_ _1959_ _1960_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__or2_2
XFILLER_116_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6221_ _3017_ vssd1 vssd1 vccd1 vccd1 _3018_ sky130_fd_sc_hd__clkbuf_2
XFILLER_104_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3208__B _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3433_ dmmu1.page_table\[0\]\[5\] dmmu1.page_table\[1\]\[5\] dmmu1.page_table\[2\]\[5\]
+ dmmu1.page_table\[3\]\[5\] _0858_ _0861_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_19_core_clock_A clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__7128__CLK clknet_leaf_29_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5704__A _2682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _2971_ dmmu0.page_table\[1\]\[12\] _2961_ vssd1 vssd1 vccd1 vccd1 _2976_ sky130_fd_sc_hd__and3_1
XFILLER_258_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _0929_ _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__nand2_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5103_ _2347_ immu_0.page_table\[13\]\[1\] _2353_ _2356_ vssd1 vssd1 vccd1 vccd1
+ _0000_ sky130_fd_sc_hd__a31o_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5423__B _2543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6083_ _2893_ _2924_ vssd1 vssd1 vccd1 vccd1 _2936_ sky130_fd_sc_hd__and2_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3295_ _0855_ _0886_ _0887_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__a21o_1
XANTENNA__4628__A1 _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3224__A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5142__C _2373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5034_ _2312_ _2302_ vssd1 vssd1 vccd1 vccd1 _2313_ sky130_fd_sc_hd__and2_1
XFILLER_272_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6985_ clknet_leaf_7_core_clock _0246_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5936_ net94 _2829_ _2846_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__a21o_1
XANTENNA__4800__A1 _2023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5867_ _2805_ dmmu1.page_table\[15\]\[8\] _2787_ _2806_ vssd1 vssd1 vccd1 vccd1 _0314_
+ sky130_fd_sc_hd__a31o_1
XFILLER_139_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3894__A _1407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6270__A _2801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4818_ _2166_ immu_1.page_table\[2\]\[5\] _2174_ vssd1 vssd1 vccd1 vccd1 _2180_ sky130_fd_sc_hd__and3_1
XFILLER_222_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5798_ _2681_ vssd1 vssd1 vccd1 vccd1 _2762_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3367__A1 _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4749_ _2137_ vssd1 vssd1 vccd1 vccd1 _2138_ sky130_fd_sc_hd__clkbuf_4
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6305__A1 _3053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7468_ net392 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_1
XFILLER_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6419_ net197 _3137_ vssd1 vssd1 vccd1 vccd1 _3138_ sky130_fd_sc_hd__and2_1
X_7399_ net338 vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4867__A1 _1981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5614__A _2370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6429__B _3137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5333__B _2497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput103 c0_sr_bus_data_o[8] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_4
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput114 c1_o_instr_long_addr[4] vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_2
XFILLER_248_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput125 c1_o_mem_addr[1] vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_2
Xinput136 c1_o_mem_data[11] vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_2
XFILLER_76_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput147 c1_o_mem_data[7] vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_2
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6084__A3 _2922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput158 c1_o_mem_long_mode vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_2
Xinput169 c1_o_req_addr[14] vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4095__A2 _1600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6445__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_21_core_clock_A clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input210_A c1_sr_bus_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3788__B _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input308_A ic0_mem_data[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5595__A2 _2632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6795__CLK clknet_leaf_80_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3358__A1 dmmu0.page_table\[1\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4412__B _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3309__A _0901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3743__S _0847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5524__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4858__A1 _1972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6339__B _3079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output527_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5897__C _2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5035__A1 _2301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6770_ clknet_leaf_90_core_clock _0031_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[9\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5586__A2 _2632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3982_ _1456_ _1494_ _1441_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__o21a_1
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_3_core_clock clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_210_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5721_ _1579_ net379 net325 vssd1 vssd1 vccd1 vccd1 _2717_ sky130_fd_sc_hd__a21bo_1
XFILLER_250_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5652_ _2666_ dmmu0.page_table\[11\]\[5\] _2671_ vssd1 vssd1 vccd1 vccd1 _2677_ sky130_fd_sc_hd__and3_1
XFILLER_175_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4603_ _2046_ vssd1 vssd1 vccd1 vccd1 _2047_ sky130_fd_sc_hd__clkbuf_4
X_5583_ _2473_ dmmu0.page_table\[12\]\[2\] _2634_ vssd1 vssd1 vccd1 vccd1 _2637_ sky130_fd_sc_hd__and3_1
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3219__A _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4534_ _1999_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__buf_4
XANTENNA__6518__CLK clknet_leaf_43_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4465_ _1946_ _1931_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__and2_1
X_7253_ clknet_leaf_20_core_clock _0514_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3653__S _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5434__A _1929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3416_ _0887_ _0998_ _1000_ _1002_ _1004_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__a32o_2
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6204_ _2994_ dmmu1.page_table\[7\]\[5\] _3000_ _3008_ vssd1 vssd1 vccd1 vccd1 _0449_
+ sky130_fd_sc_hd__a31o_1
X_7184_ clknet_leaf_28_core_clock _0445_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4396_ _1895_ vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_1
XFILLER_258_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _2845_ dmmu0.page_table\[1\]\[4\] _2962_ vssd1 vssd1 vccd1 vccd1 _2967_ sky130_fd_sc_hd__and3_1
X_3347_ dmmu1.page_table\[6\]\[1\] dmmu1.page_table\[7\]\[1\] _0858_ vssd1 vssd1 vccd1
+ vccd1 _0939_ sky130_fd_sc_hd__mux2_1
XFILLER_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6668__CLK clknet_leaf_5_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6066__A3 _2922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6066_ _2914_ dmmu1.page_table\[10\]\[1\] _2922_ _2926_ vssd1 vssd1 vccd1 vccd1 _0393_
+ sky130_fd_sc_hd__a31o_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ net122 vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__inv_2
XFILLER_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3889__A _1404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _2301_ immu_0.page_table\[15\]\[1\] _2298_ _2303_ vssd1 vssd1 vccd1 vccd1
+ _0776_ sky130_fd_sc_hd__a31o_1
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6968_ clknet_leaf_90_core_clock _0229_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4234__C1 _1479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5919_ _2229_ _2830_ _2837_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__a21o_1
XFILLER_179_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_87_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6899_ clknet_leaf_76_core_clock _0160_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5328__B _2388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4001__A2 _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3563__S _1146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5344__A _1942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input160_A c1_o_mem_sel[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input258_A dcache_wb_o_dat[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5063__B _2322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input21_A c0_o_mem_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5265__A1 _2249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3799__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4394__S _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6175__A _2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5017__A1 _2301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5519__A _1925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5238__B _2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3426__S1 _0902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput407 net407 vssd1 vssd1 vccd1 vccd1 c0_i_core_int_sreg[0] sky130_fd_sc_hd__buf_2
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput418 net418 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[15] sky130_fd_sc_hd__buf_2
Xoutput429 net429 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[0] sky130_fd_sc_hd__buf_2
XANTENNA__3473__S _0881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5254__A _2447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4250_ net114 immu_1.high_addr_off\[4\] vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__nand2_1
XFILLER_234_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6069__B _2924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3201_ net221 _0819_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__and2_1
X_4181_ immu_1.page_table\[2\]\[7\] immu_1.page_table\[3\]\[7\] _1493_ vssd1 vssd1
+ vccd1 vccd1 _1688_ sky130_fd_sc_hd__mux2_1
XFILLER_234_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6085__A _2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_255_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6822_ clknet_leaf_59_core_clock _0083_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4216__C1 _1432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6753_ clknet_leaf_88_core_clock _0014_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3965_ _1423_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3648__S _1169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5429__A _2312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5704_ _2682_ dmmu0.page_table\[2\]\[5\] _2702_ vssd1 vssd1 vccd1 vccd1 _2708_ sky130_fd_sc_hd__and3_1
XANTENNA__4333__A _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6684_ clknet_leaf_42_core_clock _0754_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3896_ net385 net2 net3 vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__nor3b_4
XANTENNA__3990__A1 _1419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5635_ _2370_ vssd1 vssd1 vccd1 vccd1 _2666_ sky130_fd_sc_hd__clkbuf_4
XFILLER_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5566_ _2226_ _2627_ _2630_ immu_0.page_table\[0\]\[2\] vssd1 vssd1 vccd1 vccd1 _0189_
+ sky130_fd_sc_hd__o22a_1
XFILLER_275_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7305_ clknet_leaf_3_core_clock _0566_ vssd1 vssd1 vccd1 vccd1 dmmu1.long_off_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4517_ net209 vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__buf_4
X_5497_ net97 _2593_ vssd1 vssd1 vccd1 vccd1 _2595_ sky130_fd_sc_hd__and2_1
XANTENNA__5164__A _2384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7236_ clknet_leaf_24_core_clock _0497_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4448_ net98 vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__clkbuf_8
XFILLER_278_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4298__A2 _1796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4379_ net117 immu_1.high_addr_off\[7\] vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__xor2_1
XFILLER_98_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7167_ clknet_leaf_4_core_clock _0428_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_258_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6118_ _2948_ dmmu1.page_table\[9\]\[10\] _2941_ _2956_ vssd1 vssd1 vccd1 vccd1 _0415_
+ sky130_fd_sc_hd__a31o_1
XFILLER_246_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6039__A3 _2902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7098_ clknet_leaf_35_core_clock _0359_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5247__A1 _2224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6049_ _2893_ _2904_ vssd1 vssd1 vccd1 vccd1 _2915_ sky130_fd_sc_hd__and2_1
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4508__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3353__S0 _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6211__A3 _3000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5339__A _1937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3408__S1 _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6833__CLK clknet_leaf_66_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input375_A ic1_wb_adr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4525__A3 _1963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5722__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3733__A1 _0868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input69_A c0_o_req_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4389__S _0811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5074__A _1928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4289__A2 _1791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5521__B _2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3249__A0 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4418__A _1373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5789__A2 _2748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3322__A _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5948__S _2848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6202__A3 _3000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6352__B _2170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5410__A1 _2531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4153__A _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3750_ net145 net40 _1322_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__mux2_2
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3681_ _0868_ _1262_ _0872_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7464__A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5420_ _2546_ immu_0.page_table\[6\]\[4\] _2541_ _2548_ vssd1 vssd1 vccd1 vccd1 _0125_
+ sky130_fd_sc_hd__a31o_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4516__A3 _1964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4072__S1 _1581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5351_ _2503_ immu_0.page_table\[9\]\[9\] _2495_ _2507_ vssd1 vssd1 vccd1 vccd1 _0097_
+ sky130_fd_sc_hd__a31o_1
XFILLER_114_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4302_ net115 immu_1.high_addr_off\[5\] vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__or2_1
X_5282_ _2230_ _2462_ _2468_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__a21o_1
XFILLER_114_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6269__A3 _3038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5477__A1 _2576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4233_ _1424_ _1738_ vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__or2_1
X_7021_ clknet_leaf_82_core_clock _0282_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3216__B _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4164_ _1516_ _1665_ _1667_ _1671_ _1553_ vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__a311o_1
XFILLER_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5431__B _2543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4095_ _1479_ _1600_ _1603_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__a21o_1
XANTENNA__4328__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3232__A _0837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6805_ clknet_leaf_82_core_clock _0066_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_223_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6262__B _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4997_ _2284_ immu_1.page_table\[15\]\[6\] _2282_ vssd1 vssd1 vccd1 vccd1 _2290_
+ sky130_fd_sc_hd__and3_1
XFILLER_210_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5401__A1 _2531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6856__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6736_ clknet_leaf_66_core_clock _0806_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[12\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3948_ net385 net107 net108 vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__or3b_4
XFILLER_211_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3963__A1 _1416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6667_ clknet_leaf_9_core_clock _0737_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3879_ net252 _1397_ _1386_ vssd1 vssd1 vccd1 vccd1 _1398_ sky130_fd_sc_hd__mux2_4
X_5618_ _2230_ _2650_ _2657_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__a21o_1
XFILLER_164_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4507__A3 _1964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6598_ clknet_leaf_56_core_clock _0668_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4063__S1 _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5606__B _2296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3715__A1 _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5549_ _2223_ _2623_ _2625_ immu_0.page_table\[1\]\[1\] vssd1 vssd1 vccd1 vccd1 _0177_
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7219_ clknet_leaf_27_core_clock _0480_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[5\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6437__B _3137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5341__B _2497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input123_A c1_o_mem_addr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3326__S0 _0897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6432__A3 _3135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6453__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5069__A _1922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4701__A _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3317__A _0900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7161__CLK clknet_leaf_9_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5532__A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6729__CLK clknet_leaf_66_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3890__A0 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3987__A _1499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5678__S _2690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7459__A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6363__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6879__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4920_ _2237_ dmmu0.page_table\[0\]\[8\] _2221_ vssd1 vssd1 vccd1 vccd1 _2246_ sky130_fd_sc_hd__and3_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_42_core_clock clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_221_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4851_ _2084_ _2193_ vssd1 vssd1 vccd1 vccd1 _2196_ sky130_fd_sc_hd__or2_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4198__A1 _1553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3802_ _1352_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_1
XFILLER_60_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4782_ _2150_ immu_1.page_table\[4\]\[1\] _2157_ vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__and3_1
XFILLER_20_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6521_ clknet_leaf_43_core_clock _0591_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3733_ _0868_ _1311_ _1313_ _0854_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__o211a_1
XFILLER_186_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5707__A _2709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6452_ _3153_ _0809_ _0810_ net213 net212 vssd1 vssd1 vccd1 vccd1 _3155_ sky130_fd_sc_hd__a311o_1
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3664_ _0909_ _1243_ _1245_ _0905_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__o211a_1
XFILLER_134_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5403_ _2531_ immu_0.page_table\[7\]\[9\] _2525_ _2537_ vssd1 vssd1 vccd1 vccd1 _0119_
+ sky130_fd_sc_hd__a31o_1
XFILLER_146_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6383_ _3114_ vssd1 vssd1 vccd1 vccd1 _3115_ sky130_fd_sc_hd__clkbuf_2
X_3595_ dmmu0.page_table\[4\]\[9\] dmmu0.page_table\[5\]\[9\] _1169_ vssd1 vssd1 vccd1
+ vccd1 _1179_ sky130_fd_sc_hd__mux2_1
XANTENNA__3227__A _0834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5334_ _2489_ immu_0.page_table\[9\]\[1\] _2495_ _2498_ vssd1 vssd1 vccd1 vccd1 _0089_
+ sky130_fd_sc_hd__a31o_1
XFILLER_125_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5265_ _2249_ _2441_ _2457_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__a21o_1
XFILLER_248_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3661__S _0896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4984__C _2282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5442__A _2561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7004_ clknet_leaf_36_core_clock _0265_ vssd1 vssd1 vccd1 vccd1 immu_1.high_addr_off\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4216_ _1423_ _1720_ _1722_ _1432_ vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__o211a_1
XANTENNA__4122__B2 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5196_ _2400_ dmmu0.page_table\[8\]\[1\] _2411_ vssd1 vssd1 vccd1 vccd1 _2413_ sky130_fd_sc_hd__and3_1
XFILLER_68_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6257__B _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4673__A2 _2083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_81_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_core_clock
+ sky130_fd_sc_hd__clkbuf_16
X_4147_ immu_1.page_table\[12\]\[6\] immu_1.page_table\[13\]\[6\] _1453_ vssd1 vssd1
+ vccd1 vccd1 _1655_ sky130_fd_sc_hd__mux2_1
XANTENNA__3881__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4078_ _1530_ _1582_ _1587_ _1457_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__a211oi_4
XANTENNA__5622__A1 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3897__A _1410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_core_clock_A clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5925__A2 _2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7034__CLK clknet_leaf_13_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6719_ clknet_leaf_63_core_clock _0789_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5617__A _2655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4521__A _1989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7184__CLK clknet_leaf_28_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6448__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput590 net590 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[13] sky130_fd_sc_hd__buf_2
XFILLER_160_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5352__A _2314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input240_A dcache_wb_adr[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input338_A ic1_mem_data[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6167__B _2983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5861__A1 _2618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3872__A0 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5613__A1 _2224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3746__S _1322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3973__C _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output557_A net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3380_ _0921_ _0970_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__and2_1
XFILLER_69_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6358__A _1910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5262__A _2447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5050_ _2316_ immu_0.page_table\[14\]\[2\] _2320_ _2324_ vssd1 vssd1 vccd1 vccd1
+ _0788_ sky130_fd_sc_hd__a31o_1
XANTENNA__4104__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6077__B _2924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4001_ _1424_ _1510_ _1512_ net315 vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__o211a_1
XANTENNA__5852__A1 _2618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3863__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4606__A _2038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5952_ dmmu0.long_off_reg\[6\] _1942_ _2848_ vssd1 vssd1 vccd1 vccd1 _2855_ sky130_fd_sc_hd__mux2_1
XFILLER_213_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4903_ _2232_ vssd1 vssd1 vccd1 vccd1 _2233_ sky130_fd_sc_hd__buf_4
X_5883_ _2223_ _2812_ _2816_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__a21o_1
XFILLER_33_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4834_ _1896_ vssd1 vssd1 vccd1 vccd1 _2190_ sky130_fd_sc_hd__buf_4
XFILLER_166_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4040__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4765_ _2016_ _2138_ _2147_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__a21o_1
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5383__A3 _2525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6504_ clknet_leaf_59_core_clock _0574_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3716_ _0905_ _1292_ _1296_ net18 vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__a211o_1
X_7484_ net166 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__buf_2
X_4696_ _2105_ vssd1 vssd1 vccd1 vccd1 _2106_ sky130_fd_sc_hd__buf_2
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6435_ net208 _3137_ vssd1 vssd1 vccd1 vccd1 _3146_ sky130_fd_sc_hd__and2_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3647_ _1229_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_1
XFILLER_146_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6366_ _3101_ dmmu1.page_table\[2\]\[5\] _3096_ _3105_ vssd1 vssd1 vccd1 vccd1 _0514_
+ sky130_fd_sc_hd__a31o_1
XFILLER_283_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3578_ _1155_ _1157_ _0874_ _1161_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__o211a_2
XFILLER_283_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5317_ _1942_ _2482_ vssd1 vssd1 vccd1 vccd1 _2488_ sky130_fd_sc_hd__and2_1
XFILLER_114_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6268__A _2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6297_ _3053_ dmmu1.page_table\[4\]\[3\] _3058_ _3064_ vssd1 vssd1 vccd1 vccd1 _0486_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__5172__A _2384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput307 ic0_mem_data[8] vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3529__S0 _0891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput318 ic0_wb_adr[3] vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_2
Xinput329 ic0_wb_we vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__buf_2
X_5248_ _2447_ dmmu0.page_table\[7\]\[2\] _2445_ vssd1 vssd1 vccd1 vccd1 _2449_ sky130_fd_sc_hd__and3_1
XFILLER_248_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5843__A1 _2618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5179_ _2400_ dmmu0.page_table\[9\]\[8\] _2392_ vssd1 vssd1 vccd1 vccd1 _2402_ sky130_fd_sc_hd__and3_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3777__D _1279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3385__A2 _0929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input190_A c1_sr_bus_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input288_A ic0_mem_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6574__CLK clknet_leaf_46_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5066__B _2322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input51_A c0_o_mem_high_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5082__A _1940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6917__CLK clknet_leaf_58_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4022__A0 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output674_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3476__S _0881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4799__C _2157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4550_ _1977_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__buf_6
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3501_ _0874_ _1082_ _1086_ _1034_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__a211o_2
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4481_ net190 net189 vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__nand2_1
XFILLER_128_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6220_ _2919_ _2118_ vssd1 vssd1 vccd1 vccd1 _3017_ sky130_fd_sc_hd__or2_1
X_3432_ _0993_ _1006_ _1007_ _1020_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__o31a_4
XFILLER_143_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _0921_ _0947_ _0954_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__o21ai_1
X_6151_ net94 _2959_ _2975_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__a21o_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6078__A1 _2932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3505__A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5102_ _1928_ _2355_ vssd1 vssd1 vccd1 vccd1 _2356_ sky130_fd_sc_hd__and2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ net123 vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__buf_4
X_6082_ _2932_ dmmu1.page_table\[10\]\[8\] _2922_ _2935_ vssd1 vssd1 vccd1 vccd1 _0400_
+ sky130_fd_sc_hd__a31o_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5825__A1 _2242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3224__B _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ net104 vssd1 vssd1 vccd1 vccd1 _2312_ sky130_fd_sc_hd__buf_4
XFILLER_285_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6984_ clknet_leaf_7_core_clock _0245_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5935_ _2845_ dmmu0.page_table\[5\]\[11\] _2831_ vssd1 vssd1 vccd1 vccd1 _2846_ sky130_fd_sc_hd__and3_1
XFILLER_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4800__A2 _2155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5866_ _1985_ _2789_ vssd1 vssd1 vccd1 vccd1 _2806_ sky130_fd_sc_hd__and2_1
XANTENNA__6002__A1 _2884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6597__CLK clknet_leaf_53_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4817_ _2012_ _2172_ _2179_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__a21o_1
XANTENNA__6270__B _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5797_ _1948_ _2748_ _2761_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__a21o_1
XFILLER_166_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4071__A _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4748_ _2000_ _2136_ vssd1 vssd1 vccd1 vccd1 _2137_ sky130_fd_sc_hd__nor2_1
XFILLER_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7467_ net391 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__clkbuf_1
XFILLER_162_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4679_ _2016_ _2083_ _2094_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__a21o_1
XFILLER_208_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7382__A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6418_ _3136_ vssd1 vssd1 vccd1 vccd1 _3137_ sky130_fd_sc_hd__buf_2
X_7398_ net337 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_1
XFILLER_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4867__A2 _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6349_ _2919_ _2170_ vssd1 vssd1 vccd1 vccd1 _3094_ sky130_fd_sc_hd__or2_1
XFILLER_115_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput104 c0_sr_bus_data_o[9] vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_4
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput115 c1_o_instr_long_addr[5] vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5816__A1 _2229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput126 c1_o_mem_addr[2] vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_2
Xinput137 c1_o_mem_data[12] vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_2
Xinput148 c1_o_mem_data[8] vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_2
XFILLER_88_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput159 c1_o_mem_req vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_1
XFILLER_248_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6445__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4246__A _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6241__A1 _3026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input203_A c1_sr_bus_data_o[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input99_A c0_sr_bus_data_o[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5347__A3 _2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4555__A1 _2014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5805__A _2216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4858__A2 _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3325__A _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5243__C _2445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3818__A0 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6480__A1 inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6232__A1 _3010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3981_ immu_1.page_table\[0\]\[1\] immu_1.page_table\[1\]\[1\] immu_1.page_table\[8\]\[1\]
+ immu_1.page_table\[9\]\[1\] _1493_ net369 vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__mux4_2
XANTENNA__5686__S _2690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7467__A net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5720_ _2253_ _2699_ _2716_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__a21o_1
XANTENNA__6371__A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5651_ _2233_ _2669_ _2676_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__a21o_1
XFILLER_148_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5338__A3 _2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4602_ _2000_ _2045_ vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__nor2_1
XANTENNA__4546__A1 _2008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5582_ _2224_ _2632_ _2636_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__a21o_1
XFILLER_190_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4533_ _1998_ vssd1 vssd1 vccd1 vccd1 _1999_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__6299__A1 _3053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5715__A _2709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7252_ clknet_leaf_24_core_clock _0513_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4464_ net103 vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__buf_6
XANTENNA__7245__CLK clknet_leaf_26_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5434__B _2555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6203_ _2799_ _3002_ vssd1 vssd1 vccd1 vccd1 _3008_ sky130_fd_sc_hd__and2_1
X_3415_ _0881_ _1003_ _0874_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__o21a_1
X_7183_ clknet_leaf_15_core_clock _0444_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4395_ net273 _1894_ _0811_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__mux2_4
XANTENNA__5510__A3 _2591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3235__A _0839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _2229_ _2960_ _2966_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__a21o_1
X_3346_ _0881_ _0937_ _0887_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__a21o_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6065_ _2791_ _2924_ vssd1 vssd1 vccd1 vccd1 _2926_ sky130_fd_sc_hd__and2_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3277_ dmmu1.page_table\[10\]\[0\] dmmu1.page_table\[11\]\[0\] _0858_ vssd1 vssd1
+ vccd1 vccd1 _0870_ sky130_fd_sc_hd__mux2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6471__A1 _1981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _1928_ _2302_ vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__and2_1
XFILLER_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4066__A net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ clknet_leaf_89_core_clock _0228_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_214_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6281__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5918_ _2834_ dmmu0.page_table\[5\]\[3\] _2832_ vssd1 vssd1 vccd1 vccd1 _2837_ sky130_fd_sc_hd__and3_1
XANTENNA__4785__A1 _2008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6898_ clknet_leaf_76_core_clock _0159_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5849_ _2618_ dmmu1.page_table\[15\]\[2\] _2787_ _2794_ vssd1 vssd1 vccd1 vccd1 _0308_
+ sky130_fd_sc_hd__a31o_1
XFILLER_21_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5625__A _2655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5344__B _2497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6612__CLK clknet_leaf_54_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input153_A c1_o_mem_high_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6456__A _2084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input320_A ic0_wb_adr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3799__B _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6175__B _2983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input14_A c0_o_mem_addr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5017__A2 immu_0.page_table\[15\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6191__A _1968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3984__C1 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4528__A1 _1976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3754__S _1322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput408 net408 vssd1 vssd1 vccd1 vccd1 c0_i_core_int_sreg[1] sky130_fd_sc_hd__buf_2
XFILLER_172_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput419 net419 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[1] sky130_fd_sc_hd__buf_2
XFILLER_99_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output637_A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3200_ _0820_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4700__A1 _2008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4180_ _1676_ _1685_ _1682_ net107 vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__o31ai_1
XFILLER_95_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6821_ clknet_leaf_61_core_clock _0082_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_250_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4614__A _1897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6752_ clknet_leaf_86_core_clock _0013_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4767__A1 _2019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3964_ _1471_ _1476_ _1410_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__or3b_2
XFILLER_50_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5429__B _2543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5703_ _2233_ _2700_ _2707_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__a21o_1
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6683_ clknet_leaf_40_core_clock _0753_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3895_ _1408_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__buf_6
XFILLER_176_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4519__A1 _1976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5148__C _2373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5634_ _2251_ _2649_ _2665_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__a21o_1
XFILLER_136_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5565_ _2223_ _2627_ _2630_ immu_0.page_table\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 _0188_
+ sky130_fd_sc_hd__o22a_1
XFILLER_163_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4987__C _2282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5445__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7304_ clknet_leaf_3_core_clock _0565_ vssd1 vssd1 vccd1 vccd1 dmmu1.long_off_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4516_ _1976_ dmmu1.page_table\[14\]\[8\] _1964_ _1986_ vssd1 vssd1 vccd1 vccd1 _0592_
+ sky130_fd_sc_hd__a31o_1
XFILLER_144_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5496_ _2588_ immu_0.page_table\[3\]\[1\] _2591_ _2594_ vssd1 vssd1 vccd1 vccd1 _0155_
+ sky130_fd_sc_hd__a31o_1
XFILLER_117_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7235_ clknet_leaf_21_core_clock _0496_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4447_ _1911_ immu_0.page_table\[11\]\[2\] _1924_ _1934_ vssd1 vssd1 vccd1 vccd1
+ _0575_ sky130_fd_sc_hd__a31o_1
XFILLER_171_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7166_ clknet_leaf_17_core_clock _0427_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6785__CLK clknet_leaf_0_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4378_ net664 _1855_ _1880_ _1881_ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__a31o_4
X_6117_ _2895_ _2943_ vssd1 vssd1 vccd1 vccd1 _2956_ sky130_fd_sc_hd__and2_1
XFILLER_219_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input6_A c0_o_instr_long_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6276__A _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3329_ _0918_ _0919_ _0921_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__a21o_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7097_ clknet_leaf_36_core_clock _0358_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6444__A1 _1898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5247__A2 _2442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _2561_ vssd1 vssd1 vccd1 vccd1 _2914_ sky130_fd_sc_hd__buf_4
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3353__S1 _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4524__A _1991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5339__B _2497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5970__A3 _2859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3574__S _0857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input270_A dcache_wb_o_dat[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4930__A1 _2251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input368_A ic1_wb_adr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5074__B _2338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_33_core_clock_A clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_150_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6186__A _1993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5090__A _2300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_32_core_clock clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7090__CLK clknet_leaf_2_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3421__A1 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6658__CLK clknet_leaf_43_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3680_ dmmu1.page_table\[10\]\[11\] dmmu1.page_table\[11\]\[11\] _0856_ vssd1 vssd1
+ vccd1 vccd1 _1262_ sky130_fd_sc_hd__mux2_1
XFILLER_145_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5350_ _2312_ _2497_ vssd1 vssd1 vccd1 vccd1 _2507_ sky130_fd_sc_hd__and2_1
XANTENNA__4921__A1 _2245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4301_ net115 immu_1.high_addr_off\[5\] vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__and2_1
XFILLER_245_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5281_ _2458_ dmmu0.page_table\[14\]\[3\] _2464_ vssd1 vssd1 vccd1 vccd1 _2468_ sky130_fd_sc_hd__and3_1
XFILLER_153_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7020_ clknet_leaf_84_core_clock _0281_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4232_ immu_0.page_table\[6\]\[8\] immu_0.page_table\[7\]\[8\] _1408_ vssd1 vssd1
+ vccd1 vccd1 _1738_ sky130_fd_sc_hd__mux2_1
XFILLER_4_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_71_core_clock clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4163_ _1581_ _1668_ _1670_ _1451_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__o211a_1
XANTENNA__6096__A _2879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6426__A1 _3128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4094_ _1535_ _1602_ _1413_ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__a21o_1
XFILLER_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4988__A1 _1967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3660__A1 _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6804_ clknet_leaf_84_core_clock _0065_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4344__A _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4996_ _1979_ _2280_ _2289_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__a21o_1
XFILLER_223_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6735_ clknet_leaf_67_core_clock _0805_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[12\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3947_ _1459_ _1460_ _1450_ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__mux2_1
XFILLER_210_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3963__A2 _1473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6666_ clknet_leaf_8_core_clock _0736_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3878_ net322 net376 _1390_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__mux2_1
XFILLER_128_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5617_ _2655_ dmmu0.page_table\[15\]\[3\] _2652_ vssd1 vssd1 vccd1 vccd1 _2657_ sky130_fd_sc_hd__and3_1
XANTENNA__5165__A1 _2224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6597_ clknet_leaf_53_core_clock _0667_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5548_ _2210_ _2623_ _2625_ immu_0.page_table\[1\]\[0\] vssd1 vssd1 vccd1 vccd1 _0176_
+ sky130_fd_sc_hd__o22a_1
XFILLER_191_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5479_ _2576_ immu_0.page_table\[4\]\[6\] _2574_ _2583_ vssd1 vssd1 vccd1 vccd1 _0149_
+ sky130_fd_sc_hd__a31o_1
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7390__A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5903__A _2819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7218_ clknet_leaf_28_core_clock _0479_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[5\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7149_ clknet_leaf_14_core_clock _0410_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3423__A _0906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3326__S1 _0902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input116_A c1_o_instr_long_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__A1 _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6196__A3 _3000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5069__B _2334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3403__A1 _0980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input81_A c0_sr_bus_addr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5156__A1 _2253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6950__CLK clknet_leaf_81_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5813__A _2762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4116__C1 _1553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3333__A net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3890__A1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6363__B _3098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4850_ _2194_ vssd1 vssd1 vccd1 vccd1 _2195_ sky130_fd_sc_hd__clkbuf_4
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6187__A3 _2980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3801_ net229 _1348_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__and2_1
XANTENNA__5395__A1 _2531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4781_ _1996_ _2155_ _2158_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__a21o_1
X_6520_ clknet_leaf_43_core_clock _0590_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3732_ net121 _1312_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__or2_1
XFILLER_158_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6451_ _3153_ mem_dcache_arb.select _0817_ _3154_ vssd1 vssd1 vccd1 vccd1 _0550_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__5147__A1 _2245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3663_ _0901_ _1244_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__or2_1
X_5402_ _2312_ _2527_ vssd1 vssd1 vccd1 vccd1 _2537_ sky130_fd_sc_hd__and2_1
XFILLER_161_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6382_ _2919_ _2187_ vssd1 vssd1 vccd1 vccd1 _3114_ sky130_fd_sc_hd__or2_1
XFILLER_133_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3594_ _1171_ _1173_ _1175_ _1177_ _0921_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__a221o_1
XFILLER_161_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5333_ _1928_ _2497_ vssd1 vssd1 vccd1 vccd1 _2498_ sky130_fd_sc_hd__and2_1
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5264_ _2447_ dmmu0.page_table\[7\]\[10\] _2444_ vssd1 vssd1 vccd1 vccd1 _2457_ sky130_fd_sc_hd__and3_1
XFILLER_125_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7003_ clknet_leaf_36_core_clock _0264_ vssd1 vssd1 vccd1 vccd1 immu_1.high_addr_off\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4215_ net313 _1721_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__or2_1
XFILLER_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5195_ _2211_ _2409_ _2412_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__a21o_1
XANTENNA__3243__A _0844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4146_ _1411_ _1641_ _1647_ _1653_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__a31o_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3881__A1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _1496_ _1583_ _1586_ _1516_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__o211a_1
XFILLER_243_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5622__A2 _2650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3633__A1 dmmu0.page_table\[9\]\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3389__S _0855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6178__A3 _2981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5386__A1 _2517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6973__CLK clknet_leaf_0_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4979_ _1960_ _2063_ vssd1 vssd1 vccd1 vccd1 _2278_ sky130_fd_sc_hd__or2_2
XANTENNA__7385__A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6718_ clknet_leaf_62_core_clock _0788_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6649_ clknet_leaf_40_core_clock _0719_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4521__B _1970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4013__S _1524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5633__A _2655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput580 net580 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[5] sky130_fd_sc_hd__buf_2
XANTENNA__6448__B _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput591 net591 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[14] sky130_fd_sc_hd__buf_2
XANTENNA__5352__B _2497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5310__A1 _2363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input233_A dcache_wb_adr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3872__A1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6464__A _2971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input400_A inner_wb_i_dat[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5613__A2 _2650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5377__A1 _2517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3483__S0 _0900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5246__C _2445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output452_A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3762__S _1322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5301__A1 _2253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4159__A _1584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6846__CLK clknet_leaf_69_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4000_ _1419_ _1511_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__or2_1
XFILLER_84_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3863__A1 _1385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5951_ _2854_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4902_ net99 vssd1 vssd1 vccd1 vccd1 _2232_ sky130_fd_sc_hd__buf_4
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5882_ _2777_ dmmu0.page_table\[6\]\[1\] _2814_ vssd1 vssd1 vccd1 vccd1 _2816_ sky130_fd_sc_hd__and3_1
XFILLER_206_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4833_ _2188_ vssd1 vssd1 vccd1 vccd1 _2189_ sky130_fd_sc_hd__buf_4
XFILLER_33_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4764_ _2134_ immu_1.page_table\[5\]\[6\] _2140_ vssd1 vssd1 vccd1 vccd1 _2147_ sky130_fd_sc_hd__and3_1
XANTENNA__4040__A1 _1410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3474__S0 _0858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6503_ clknet_leaf_60_core_clock _0573_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_267_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3715_ _0908_ _1293_ _1295_ _0917_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__o211a_1
XFILLER_146_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7483_ net165 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__buf_2
X_4695_ _1896_ vssd1 vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__buf_4
X_6434_ _1898_ dmmu1.page_table\[0\]\[7\] _3135_ _3145_ vssd1 vssd1 vccd1 vccd1 _0542_
+ sky130_fd_sc_hd__a31o_1
X_3646_ _1211_ _1228_ _0847_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__mux2_4
XFILLER_106_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6365_ net205 _3098_ vssd1 vssd1 vccd1 vccd1 _3105_ sky130_fd_sc_hd__and2_1
XANTENNA__5540__A1 _2618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3577_ _0859_ _1158_ _1160_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__a21o_1
XANTENNA__4995__C _2282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5453__A net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5316_ _2363_ immu_0.page_table\[10\]\[5\] _2480_ _2487_ vssd1 vssd1 vccd1 vccd1
+ _0082_ sky130_fd_sc_hd__a31o_1
XFILLER_142_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6296_ net203 _3060_ vssd1 vssd1 vccd1 vccd1 _3064_ sky130_fd_sc_hd__and2_1
XANTENNA__6268__B _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput308 ic0_mem_data[9] vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3529__S1 _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5247_ _2224_ _2442_ _2448_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__a21o_1
XANTENNA__4069__A _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput319 ic0_wb_adr[4] vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_2
XFILLER_88_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5178_ _2243_ _2390_ _2401_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__a21o_1
XFILLER_152_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4129_ immu_0.page_table\[10\]\[6\] immu_0.page_table\[11\]\[6\] _1601_ vssd1 vssd1
+ vccd1 vccd1 _1637_ sky130_fd_sc_hd__mux2_1
XFILLER_244_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7001__CLK clknet_leaf_37_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3420__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4008__S _1443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7151__CLK clknet_leaf_33_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6719__CLK clknet_leaf_63_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input183_A c1_sr_bus_addr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6323__A3 _3077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5531__A1 _2603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6869__CLK clknet_leaf_69_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5363__A _1935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input350_A ic1_mem_data[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5082__B _2338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input44_A c0_o_mem_data[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4098__A1 _1535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4707__A _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5062__A3 _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5538__A _2561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4442__A _1914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5770__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3500_ _0887_ _1085_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__and2_1
XFILLER_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4480_ net181 net188 vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__or2b_1
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6314__A3 _3057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3431_ _1010_ _1018_ _1019_ _0835_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__a211o_1
XANTENNA__5273__A _2443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6150_ _2971_ dmmu0.page_table\[1\]\[11\] _2961_ vssd1 vssd1 vccd1 vccd1 _2975_ sky130_fd_sc_hd__and3_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _0906_ _0949_ _0953_ _0899_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__a211o_1
XFILLER_97_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5704__C _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _1930_ _2351_ vssd1 vssd1 vccd1 vccd1 _2355_ sky130_fd_sc_hd__nor2_4
XFILLER_111_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6081_ _2891_ _2924_ vssd1 vssd1 vccd1 vccd1 _2935_ sky130_fd_sc_hd__and2_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ dmmu1.page_table\[4\]\[0\] dmmu1.page_table\[5\]\[0\] dmmu1.page_table\[6\]\[0\]
+ dmmu1.page_table\[7\]\[0\] _0865_ _0863_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__mux4_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5032_ _2301_ immu_0.page_table\[15\]\[8\] _2298_ _2311_ vssd1 vssd1 vccd1 vccd1
+ _0783_ sky130_fd_sc_hd__a31o_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4617__A _2054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6983_ clknet_leaf_78_core_clock _0244_ vssd1 vssd1 vccd1 vccd1 immu_0.high_addr_off\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_226_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7174__CLK clknet_leaf_35_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5934_ _2681_ vssd1 vssd1 vccd1 vccd1 _2845_ sky130_fd_sc_hd__buf_2
XFILLER_280_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5865_ _2561_ vssd1 vssd1 vccd1 vccd1 _2805_ sky130_fd_sc_hd__buf_4
XFILLER_221_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4816_ _2166_ immu_1.page_table\[2\]\[4\] _2174_ vssd1 vssd1 vccd1 vccd1 _2179_ sky130_fd_sc_hd__and3_1
X_5796_ _2749_ dmmu0.page_table\[13\]\[9\] _2751_ vssd1 vssd1 vccd1 vccd1 _2761_ sky130_fd_sc_hd__and3_1
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4747_ _2027_ _2117_ vssd1 vssd1 vccd1 vccd1 _2136_ sky130_fd_sc_hd__or2_4
XFILLER_147_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3772__A0 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7466_ net390 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_1
XFILLER_147_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4678_ _2089_ immu_1.page_table\[10\]\[6\] _2086_ vssd1 vssd1 vccd1 vccd1 _2094_
+ sky130_fd_sc_hd__and3_1
XANTENNA__6305__A3 _3058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6417_ _2784_ _2272_ vssd1 vssd1 vccd1 vccd1 _3136_ sky130_fd_sc_hd__nor2_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3629_ dmmu0.page_table\[12\]\[10\] dmmu0.page_table\[13\]\[10\] _0895_ vssd1 vssd1
+ vccd1 vccd1 _1212_ sky130_fd_sc_hd__mux2_1
X_7397_ net336 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5183__A _2400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6348_ _3085_ dmmu1.page_table\[3\]\[12\] _3076_ _3093_ vssd1 vssd1 vccd1 vccd1 _0508_
+ sky130_fd_sc_hd__a31o_1
XFILLER_227_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_38_core_clock_A clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_6279_ _3042_ dmmu1.page_table\[5\]\[10\] _3037_ _3052_ vssd1 vssd1 vccd1 vccd1 _0480_
+ sky130_fd_sc_hd__a31o_1
Xinput105 c0_sr_bus_we vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
Xinput116 c1_o_instr_long_addr[6] vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_2
XANTENNA__5911__A _2819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput127 c1_o_mem_addr[3] vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__buf_2
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput138 c1_o_mem_data[13] vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
XFILLER_88_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput149 c1_o_mem_data[9] vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_2
XFILLER_243_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4527__A _1993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3460__C1 _0918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5358__A _1930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input398_A inner_wb_i_dat[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4555__A2 _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6691__CLK clknet_leaf_39_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5504__A1 _2588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5805__B _2589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5093__A _2314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7047__CLK clknet_leaf_37_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5821__A _2762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7197__CLK clknet_leaf_28_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6480__A2 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4437__A _1926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3341__A _0863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5035__A3 _2298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3980_ _1443_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__buf_6
XFILLER_262_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_40_core_clock_A clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_50_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6371__B _3098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3451__C1 _0906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5650_ _2666_ dmmu0.page_table\[11\]\[4\] _2671_ vssd1 vssd1 vccd1 vccd1 _2676_ sky130_fd_sc_hd__and3_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4601_ net188 net181 _1960_ vssd1 vssd1 vccd1 vccd1 _2045_ sky130_fd_sc_hd__or3_2
XFILLER_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4546__A2 _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5581_ _2473_ dmmu0.page_table\[12\]\[1\] _2634_ vssd1 vssd1 vccd1 vccd1 _2636_ sky130_fd_sc_hd__and3_1
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3754__A0 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4532_ _1957_ _1997_ vssd1 vssd1 vccd1 vccd1 _1998_ sky130_fd_sc_hd__or2_2
XANTENNA__4900__A _2204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7251_ clknet_leaf_19_core_clock _0512_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4463_ _1939_ immu_0.page_table\[11\]\[7\] _1924_ _1945_ vssd1 vssd1 vccd1 vccd1
+ _0580_ sky130_fd_sc_hd__a31o_1
XFILLER_116_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6202_ _2994_ dmmu1.page_table\[7\]\[4\] _3000_ _3007_ vssd1 vssd1 vccd1 vccd1 _0448_
+ sky130_fd_sc_hd__a31o_1
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3414_ dmmu1.page_table\[4\]\[4\] dmmu1.page_table\[5\]\[4\] dmmu1.page_table\[6\]\[4\]
+ dmmu1.page_table\[7\]\[4\] _0865_ _0863_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__mux4_1
X_7182_ clknet_leaf_29_core_clock _0443_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[8\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_4394_ net327 net381 _0812_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__mux2_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _2845_ dmmu0.page_table\[1\]\[3\] _2962_ vssd1 vssd1 vccd1 vccd1 _2966_ sky130_fd_sc_hd__and3_1
X_3345_ dmmu1.page_table\[0\]\[1\] dmmu1.page_table\[1\]\[1\] dmmu1.page_table\[2\]\[1\]
+ dmmu1.page_table\[3\]\[1\] _0891_ _0860_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__mux4_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6064_ _2914_ dmmu1.page_table\[10\]\[0\] _2922_ _2925_ vssd1 vssd1 vccd1 vccd1 _0392_
+ sky130_fd_sc_hd__a31o_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _0868_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__clkbuf_8
XFILLER_218_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _1930_ _2296_ vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__nor2_4
XFILLER_85_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6471__A2 _3157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4347__A _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6564__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4967__A2_N _2274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6966_ clknet_leaf_86_core_clock _0227_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4234__A1 _1570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5917_ _2226_ _2830_ _2836_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__a21o_1
XFILLER_241_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4785__A2 _2155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6897_ clknet_leaf_75_core_clock _0158_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3397__S _0906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5848_ _2793_ _2789_ vssd1 vssd1 vccd1 vccd1 _2794_ sky130_fd_sc_hd__and2_1
XFILLER_194_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5734__A1 _1977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5779_ _2210_ _2748_ _2752_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__a21o_1
XANTENNA__4093__S0 _1601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7393__A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4810__A _2166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7449_ net63 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_1
XFILLER_174_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5641__A _2670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6447__C1 _1911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input146_A c1_o_mem_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6907__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4257__A _1581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input313_A ic0_wb_adr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_core_clock clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5017__A3 _2298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6472__A _2190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6191__B _2255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5973__A1 _2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5088__A _2310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3736__B1 _1316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput409 net409 vssd1 vssd1 vccd1 vccd1 c0_i_irq sky130_fd_sc_hd__buf_2
XANTENNA__5254__C _2445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4700__A2 _2101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output532_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_61_core_clock clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3770__S _0839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6587__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6382__A _2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6820_ clknet_leaf_68_core_clock _0081_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4216__A1 _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5964__A1 _2805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6751_ clknet_leaf_88_core_clock _0012_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3963_ _1416_ _1473_ _1475_ _1434_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__o211a_1
XFILLER_90_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4767__A2 _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5702_ _2682_ dmmu0.page_table\[2\]\[4\] _2702_ vssd1 vssd1 vccd1 vccd1 _2707_ sky130_fd_sc_hd__and3_1
X_6682_ clknet_leaf_41_core_clock _0752_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[7\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3894_ _1407_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__clkbuf_8
X_5633_ _2655_ dmmu0.page_table\[15\]\[11\] _2651_ vssd1 vssd1 vccd1 vccd1 _2665_
+ sky130_fd_sc_hd__and3_1
XANTENNA__5716__A1 _2249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4630__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5564_ _2628_ vssd1 vssd1 vccd1 vccd1 _2630_ sky130_fd_sc_hd__clkbuf_4
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4515_ _1985_ _1970_ vssd1 vssd1 vccd1 vccd1 _1986_ sky130_fd_sc_hd__and2_1
XANTENNA__5445__B _2559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7303_ clknet_leaf_3_core_clock _0564_ vssd1 vssd1 vccd1 vccd1 dmmu1.long_off_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_275_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5495_ net96 _2593_ vssd1 vssd1 vccd1 vccd1 _2594_ sky130_fd_sc_hd__and2_1
XFILLER_132_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7234_ clknet_leaf_26_core_clock _0495_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[4\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5164__C _2392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4446_ _1933_ _1931_ vssd1 vssd1 vccd1 vccd1 _1934_ sky130_fd_sc_hd__and2_1
X_7165_ clknet_leaf_10_core_clock _0426_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4377_ inner_wb_arbiter.o_sel_sig net245 vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__and2_1
XANTENNA__3680__S _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6116_ _2948_ dmmu1.page_table\[9\]\[9\] _2942_ _2955_ vssd1 vssd1 vccd1 vccd1 _0414_
+ sky130_fd_sc_hd__a31o_1
XFILLER_258_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3328_ _0920_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__buf_4
X_7096_ clknet_leaf_32_core_clock _0357_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6276__B _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4276__A2_N _1781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6047_ _2898_ dmmu1.page_table\[11\]\[8\] _2902_ _2913_ vssd1 vssd1 vccd1 vccd1 _0387_
+ sky130_fd_sc_hd__a31o_1
XFILLER_218_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ net119 net14 _0847_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__mux2_2
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7388__A net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6292__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6949_ clknet_leaf_7_core_clock _0210_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[12\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_241_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3855__S _1360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5636__A _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4391__A0 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input263_A dcache_wb_o_dat[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6132__A1 _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3590__S _1169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4694__A1 _1996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6186__B _2982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4715__A _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5946__A1 _1935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5410__A3 _2541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3709__B1 _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5546__A _2190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4921__A2 _2219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4300_ net2 _1786_ _1804_ _1411_ _1579_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__a221o_1
X_5280_ _2227_ _2462_ _2467_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__a21o_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4231_ immu_0.page_table\[4\]\[8\] immu_0.page_table\[5\]\[8\] _1601_ vssd1 vssd1
+ vccd1 vccd1 _1737_ sky130_fd_sc_hd__mux2_1
XFILLER_114_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5477__A3 _2574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6377__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4685__A1 _2023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5281__A _2458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4162_ _1447_ _1669_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__or2_1
XFILLER_228_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6096__B _2944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4093_ immu_0.page_table\[0\]\[5\] immu_0.page_table\[1\]\[5\] immu_0.page_table\[2\]\[5\]
+ immu_0.page_table\[3\]\[5\] _1601_ _1420_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__mux4_1
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4988__A2 _2280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4625__A _2054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6803_ clknet_leaf_81_core_clock _0064_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4995_ _2284_ immu_1.page_table\[15\]\[5\] _2282_ vssd1 vssd1 vccd1 vccd1 _2289_
+ sky130_fd_sc_hd__and3_1
XFILLER_211_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6602__CLK clknet_leaf_54_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5401__A3 _2525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6734_ clknet_leaf_66_core_clock _0804_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3946_ immu_1.page_table\[8\]\[0\] immu_1.page_table\[9\]\[0\] immu_1.page_table\[10\]\[0\]
+ immu_1.page_table\[11\]\[0\] _1437_ net367 vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__mux4_2
XFILLER_211_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4070__C1 _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3877_ _1396_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_1
X_6665_ clknet_leaf_9_core_clock _0735_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5616_ _2227_ _2650_ _2656_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__a21o_1
XFILLER_164_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5165__A2 _2390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6362__A1 _3101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6596_ clknet_leaf_53_core_clock _0666_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_219_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6752__CLK clknet_leaf_86_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5547_ _2624_ vssd1 vssd1 vccd1 vccd1 _2625_ sky130_fd_sc_hd__clkbuf_4
XFILLER_117_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6114__A1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5478_ net101 _2577_ vssd1 vssd1 vccd1 vccd1 _2583_ sky130_fd_sc_hd__and2_1
XFILLER_3_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7217_ clknet_leaf_28_core_clock _0478_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[5\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_4429_ net86 _1918_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__or2_1
XANTENNA__5903__B dmmu0.page_table\[6\]\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6287__A _3057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7108__CLK clknet_leaf_37_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7148_ clknet_leaf_34_core_clock _0409_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_274_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7079_ clknet_leaf_11_core_clock _0340_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[5\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7258__CLK clknet_leaf_25_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_274_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4535__A _1961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input109_A c1_o_icache_flush vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4600__A1 _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3403__A2 _0984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input380_A ic1_wb_sel[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4701__C _2103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input74_A c0_o_req_addr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5813__B dmmu0.page_table\[3\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6197__A _2793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5092__A1 _2347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6625__CLK clknet_leaf_54_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4445__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5919__A1 _2229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3800_ _1351_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_1
X_4780_ _2150_ immu_1.page_table\[4\]\[0\] _2157_ vssd1 vssd1 vccd1 vccd1 _2158_ sky130_fd_sc_hd__and3_1
XANTENNA__4052__C1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ dmmu1.page_table\[12\]\[12\] dmmu1.page_table\[13\]\[12\] net120 vssd1 vssd1
+ vccd1 vccd1 _1312_ sky130_fd_sc_hd__mux2_1
XANTENNA__6775__CLK clknet_leaf_81_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6344__A1 _3085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6450_ net710 _0809_ vssd1 vssd1 vccd1 vccd1 _3154_ sky130_fd_sc_hd__nor2_1
XANTENNA__5147__A2 _2369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3662_ dmmu0.page_table\[12\]\[11\] dmmu0.page_table\[13\]\[11\] _1169_ vssd1 vssd1
+ vccd1 vccd1 _1244_ sky130_fd_sc_hd__mux2_1
XANTENNA__5707__C _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4355__B1 _1516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5401_ _2531_ immu_0.page_table\[7\]\[8\] _2525_ _2536_ vssd1 vssd1 vccd1 vccd1 _0118_
+ sky130_fd_sc_hd__a31o_1
X_6381_ _3112_ dmmu1.page_table\[2\]\[12\] _3095_ _3113_ vssd1 vssd1 vccd1 vccd1 _0521_
+ sky130_fd_sc_hd__a31o_1
XFILLER_173_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3593_ _0908_ _1176_ _0917_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__a21oi_1
XFILLER_161_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7491__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5332_ _1930_ _2388_ vssd1 vssd1 vccd1 vccd1 _2497_ sky130_fd_sc_hd__nor2_4
XFILLER_114_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5263_ _2247_ _2442_ _2456_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__a21o_1
XANTENNA__4658__A1 _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4214_ immu_0.page_table\[12\]\[7\] immu_0.page_table\[13\]\[7\] net312 vssd1 vssd1
+ vccd1 vccd1 _1721_ sky130_fd_sc_hd__mux2_1
X_7002_ clknet_leaf_37_core_clock _0263_ vssd1 vssd1 vccd1 vccd1 immu_1.high_addr_off\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5194_ _2400_ dmmu0.page_table\[8\]\[0\] _2411_ vssd1 vssd1 vccd1 vccd1 _2412_ sky130_fd_sc_hd__and3_1
XFILLER_205_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4145_ net2 _1652_ _1360_ vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__a21o_1
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4076_ _1584_ _1585_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__or2_1
XFILLER_243_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5083__A1 _2332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4830__A1 _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4978_ _1989_ _2273_ _2277_ immu_1.page_table\[0\]\[10\] vssd1 vssd1 vccd1 vccd1
+ _0763_ sky130_fd_sc_hd__o22a_1
XFILLER_196_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6717_ clknet_leaf_63_core_clock _0787_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3929_ net366 vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__buf_6
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5617__C _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6648_ clknet_leaf_38_core_clock _0718_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3418__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6579_ clknet_leaf_49_core_clock _0649_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[10\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4897__A1 _2227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5914__A _2834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput570 net570 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[10] sky130_fd_sc_hd__buf_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput581 net581 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[6] sky130_fd_sc_hd__buf_2
XANTENNA__6448__C _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput592 net592 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[15] sky130_fd_sc_hd__buf_2
XANTENNA__7080__CLK clknet_leaf_11_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5861__A3 _2787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6648__CLK clknet_leaf_38_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input226_A dcache_mem_o_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4821__A1 _2016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6798__CLK clknet_leaf_10_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_45_core_clock_A clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_24_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3483__S1 _0902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5824__A _2777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output445_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5262__C _2445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5852__A3 _2787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5950_ dmmu0.long_off_reg\[5\] _1940_ _2848_ vssd1 vssd1 vccd1 vccd1 _2854_ sky130_fd_sc_hd__mux2_1
XFILLER_225_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4273__C1 _1553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4606__C _2049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4901_ _2230_ _2219_ _2231_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__a21o_1
XFILLER_280_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5881_ _2210_ _2812_ _2815_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__a21o_1
XFILLER_233_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4832_ _1999_ _2187_ vssd1 vssd1 vccd1 vccd1 _2188_ sky130_fd_sc_hd__or2_1
XANTENNA__4903__A _2232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4763_ _2014_ _2138_ _2146_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__a21o_1
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3474__S1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4114__S _1438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6502_ _3183_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__clkbuf_1
X_3714_ net16 _1294_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__or2_1
X_4694_ _1996_ _2101_ _2104_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__a21o_1
X_7482_ net179 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_2
XFILLER_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6433_ net207 _3137_ vssd1 vssd1 vccd1 vccd1 _3145_ sky130_fd_sc_hd__and2_1
X_3645_ _1009_ _1221_ _1227_ net53 vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__a22o_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5232__B1_N net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3576_ _0868_ _1159_ _0854_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__a21o_1
X_6364_ _3101_ dmmu1.page_table\[2\]\[4\] _3096_ _3104_ vssd1 vssd1 vccd1 vccd1 _0513_
+ sky130_fd_sc_hd__a31o_1
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5453__B _2559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5315_ _1940_ _2482_ vssd1 vssd1 vccd1 vccd1 _2487_ sky130_fd_sc_hd__and2_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6295_ _3053_ dmmu1.page_table\[4\]\[2\] _3058_ _3063_ vssd1 vssd1 vccd1 vccd1 _0485_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__3254__A _0850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5172__C _2392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput309 ic0_wb_adr[0] vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_2
X_5246_ _2447_ dmmu0.page_table\[7\]\[1\] _2445_ vssd1 vssd1 vccd1 vccd1 _2448_ sky130_fd_sc_hd__and3_1
XFILLER_275_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5843__A3 _2787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5177_ _2400_ dmmu0.page_table\[9\]\[7\] _2392_ vssd1 vssd1 vccd1 vccd1 _2401_ sky130_fd_sc_hd__and3_1
XFILLER_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4128_ _1570_ _1635_ vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__or2_2
XFILLER_244_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5056__A1 _2316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4059_ inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__buf_4
XANTENNA__4085__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4264__C1 _1553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7396__A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5909__A _2443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4016__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6308__A1 _3069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3863__S _1386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5644__A _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input176_A c1_o_req_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5363__B _2512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input343_A ic1_mem_data[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5295__A1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input37_A c0_o_mem_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4707__B immu_1.page_table\[9\]\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5819__A _2762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4442__B _1930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5770__A2 _2729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output562_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6813__CLK clknet_leaf_1_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3430_ _1009_ net19 vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__and2b_1
XFILLER_116_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6369__B _3098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5273__B _2318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3361_ _0948_ _0950_ _0952_ _0918_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__o211a_1
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5100_ _2347_ immu_0.page_table\[13\]\[0\] _2353_ _2354_ vssd1 vssd1 vccd1 vccd1
+ _0808_ sky130_fd_sc_hd__a31o_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6080_ _2932_ dmmu1.page_table\[10\]\[7\] _2922_ _2934_ vssd1 vssd1 vccd1 vccd1 _0399_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__6078__A3 _2922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _0869_ _0884_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__or2_1
XFILLER_111_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5286__A1 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _2310_ _2302_ vssd1 vssd1 vccd1 vccd1 _2311_ sky130_fd_sc_hd__and2_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6385__A _2784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3392__S0 _0858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5038__A1 _2301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6982_ clknet_leaf_78_core_clock _0243_ vssd1 vssd1 vccd1 vccd1 immu_0.high_addr_off\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_241_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5933_ _1950_ _2829_ _2844_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__a21o_1
XFILLER_241_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5864_ _2618_ dmmu1.page_table\[15\]\[7\] _2787_ _2804_ vssd1 vssd1 vccd1 vccd1 _0313_
+ sky130_fd_sc_hd__a31o_1
XFILLER_33_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4815_ _2010_ _2172_ _2178_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__a21o_1
XANTENNA__6002__A3 _2878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5210__A1 _2243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5795_ _1946_ _2748_ _2760_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__a21o_1
X_4746_ _2025_ _2119_ _2135_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__a21o_1
XFILLER_193_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7465_ net404 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_1
X_4677_ _2014_ _2083_ _2093_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__a21o_1
XFILLER_107_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5464__A _1925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6416_ _3134_ vssd1 vssd1 vccd1 vccd1 _3135_ sky130_fd_sc_hd__clkbuf_4
XFILLER_174_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3628_ _0995_ _1204_ _1210_ net158 vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__a22o_2
XFILLER_162_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7396_ net335 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5183__B dmmu0.page_table\[9\]\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6347_ net200 _3078_ vssd1 vssd1 vccd1 vccd1 _3093_ sky130_fd_sc_hd__and2_1
XFILLER_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3559_ _1088_ _1128_ _1143_ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__a21o_4
XFILLER_115_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6278_ _2895_ _3039_ vssd1 vssd1 vccd1 vccd1 _3052_ sky130_fd_sc_hd__and2_1
XFILLER_88_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput106 c1_o_c_data_page vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_2
Xinput117 c1_o_instr_long_addr[7] vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput128 c1_o_mem_addr[4] vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_2
Xinput139 c1_o_mem_data[14] vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_2
X_5229_ _2099_ _2429_ vssd1 vssd1 vccd1 vccd1 _2434_ sky130_fd_sc_hd__nor2_2
XFILLER_276_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4808__A _2166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3383__S0 _0898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5029__A1 _2301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_core_clock clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_244_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6241__A3 _3019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3858__S _1360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5358__B _2407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5201__A1 _2230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6836__CLK clknet_leaf_69_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input293_A ic0_mem_data[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5374__A _2310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5093__B _2338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6986__CLK clknet_leaf_7_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_51_core_clock clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5268__A1 _2251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3622__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3374__S0 _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output408_A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6232__A3 _3019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5440__A1 _2546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3768__S _0839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4600_ _2025_ _2029_ _2044_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__a21o_1
XFILLER_30_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5580_ _2211_ _2632_ _2635_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__a21o_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_90_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4531_ _1953_ net196 net195 vssd1 vssd1 vccd1 vccd1 _1997_ sky130_fd_sc_hd__or3b_4
XFILLER_129_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6299__A3 _3058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7250_ clknet_leaf_20_core_clock _0511_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4462_ _1944_ _1931_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__and2_1
XFILLER_264_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6201_ _2797_ _3002_ vssd1 vssd1 vccd1 vccd1 _3007_ sky130_fd_sc_hd__and2_1
XANTENNA__3516__B _1101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3506__A1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3413_ _0855_ _1001_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__or2_1
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7181_ clknet_leaf_29_core_clock _0442_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[8\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_4393_ _1893_ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__clkbuf_1
XFILLER_98_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3344_ _0872_ _0935_ _0874_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__a21o_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6132_ _2226_ _2960_ _2965_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__a21o_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__A1 _2243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3275_ net121 vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__inv_2
X_6063_ _2879_ _2924_ vssd1 vssd1 vccd1 vccd1 _2925_ sky130_fd_sc_hd__and2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7141__CLK clknet_leaf_27_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3532__A _0863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5014_ _2300_ vssd1 vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__clkbuf_4
XFILLER_285_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6709__CLK clknet_leaf_63_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7291__CLK clknet_leaf_44_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6965_ clknet_leaf_87_core_clock _0226_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3678__S _1146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5459__A _2314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5916_ _2834_ dmmu0.page_table\[5\]\[2\] _2832_ vssd1 vssd1 vccd1 vccd1 _2836_ sky130_fd_sc_hd__and3_1
X_6896_ clknet_leaf_82_core_clock _0157_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5847_ net202 vssd1 vssd1 vccd1 vccd1 _2793_ sky130_fd_sc_hd__buf_2
XFILLER_21_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5778_ _2749_ dmmu0.page_table\[13\]\[0\] _2751_ vssd1 vssd1 vccd1 vccd1 _2752_ sky130_fd_sc_hd__and3_1
XANTENNA__4093__S1 _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4729_ _2008_ _2120_ _2126_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__a21o_1
XANTENNA__5194__A _2400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3707__A _0901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5625__C _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7448_ net62 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_1
XFILLER_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5498__A1 _2588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7379_ clknet_leaf_19_core_clock vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_2
XANTENNA__5922__A _2834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3442__A _0863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input139_A c1_o_mem_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3681__B1 _0872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input306_A ic0_mem_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3588__S _1169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5422__A1 _2546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4225__A2 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3984__A1 _1487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5088__B _2338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3984__B2 _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4528__A3 _1963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7014__CLK clknet_leaf_38_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3617__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7164__CLK clknet_leaf_9_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5832__A _2777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4448__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output525_A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6382__B _2187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5413__A1 _2531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5279__A _2458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6750_ clknet_leaf_89_core_clock _0011_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4183__A _1442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3962_ _1467_ _1474_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__or2_1
XFILLER_250_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5701_ _2230_ _2700_ _2706_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__a21o_1
X_6681_ clknet_leaf_41_core_clock _0751_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[7\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3893_ net312 vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__buf_6
XFILLER_231_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7494__A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5632_ _2249_ _2649_ _2664_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__a21o_1
XANTENNA__4911__A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4519__A3 _1964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4630__B net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5563_ _1926_ _2627_ _2629_ immu_0.page_table\[0\]\[0\] vssd1 vssd1 vccd1 vccd1 _0187_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_191_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7302_ clknet_leaf_62_core_clock _0563_ vssd1 vssd1 vccd1 vccd1 inner_wb_arbiter.o_sel_sig
+ sky130_fd_sc_hd__dfxtp_4
X_4514_ net208 vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__buf_4
XFILLER_191_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5494_ _1922_ _2589_ vssd1 vssd1 vccd1 vccd1 _2593_ sky130_fd_sc_hd__nor2_4
XFILLER_117_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7233_ clknet_leaf_26_core_clock _0494_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[4\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_278_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4445_ net97 vssd1 vssd1 vccd1 vccd1 _1933_ sky130_fd_sc_hd__buf_6
XANTENNA__3961__S _1407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4225__B1_N _1731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5742__A _2216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4152__A1 immu_1.page_table\[9\]\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7164_ clknet_leaf_9_core_clock _0425_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6531__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4376_ _1441_ _1864_ _1873_ _1879_ _0813_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__a311o_2
X_6115_ _2893_ _2944_ vssd1 vssd1 vccd1 vccd1 _2955_ sky130_fd_sc_hd__and2_1
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3327_ net18 vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__inv_2
XFILLER_86_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7095_ clknet_leaf_37_core_clock _0356_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_258_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3262__A _0854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6444__A3 _3134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6046_ _2891_ _2904_ vssd1 vssd1 vccd1 vccd1 _2913_ sky130_fd_sc_hd__and2_1
XFILLER_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3258_ _0852_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_2
XFILLER_224_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6681__CLK clknet_leaf_41_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3189_ icache_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__buf_6
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6292__B _3060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3415__B1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6948_ clknet_leaf_81_core_clock _0209_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[12\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7037__CLK clknet_leaf_12_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3510__S0 _0897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6879_ clknet_leaf_71_core_clock _0140_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[5\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3718__A1 _0957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7187__CLK clknet_leaf_28_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4032__S _1472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6132__A2 _2960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5652__A _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input256_A dcache_wb_o_dat[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_core_clock clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4694__A2 _2101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4268__A _1442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5643__A1 _2211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5099__A _1926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3709__A1 _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6554__CLK clknet_leaf_50_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4230_ _1734_ _1735_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__xnor2_2
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4685__A2 _2083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3342__C1 _0854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4161_ immu_1.page_table\[2\]\[6\] immu_1.page_table\[3\]\[6\] _1437_ vssd1 vssd1
+ vccd1 vccd1 _1669_ sky130_fd_sc_hd__mux2_1
XFILLER_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4092_ _1408_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__buf_6
XANTENNA__6426__A3 _3135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5634__A1 _2251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7489__A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_255_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4906__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6802_ clknet_leaf_6_core_clock _0063_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[7\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4117__S _1448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4994_ _1977_ _2280_ _2288_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__a21o_1
XFILLER_251_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6733_ clknet_leaf_63_core_clock _0803_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3945_ immu_1.page_table\[12\]\[0\] immu_1.page_table\[13\]\[0\] immu_1.page_table\[14\]\[0\]
+ immu_1.page_table\[15\]\[0\] _1437_ net367 vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__mux4_1
XFILLER_149_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6664_ clknet_leaf_8_core_clock _0734_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3876_ net251 _1395_ _1386_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__mux2_4
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5615_ _2655_ dmmu0.page_table\[15\]\[2\] _2652_ vssd1 vssd1 vccd1 vccd1 _2656_ sky130_fd_sc_hd__and3_1
XFILLER_176_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6595_ clknet_leaf_59_core_clock _0665_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_117_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5546_ _2190_ _2622_ vssd1 vssd1 vccd1 vccd1 _2624_ sky130_fd_sc_hd__nand2_1
XFILLER_129_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3691__S _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5477_ _2576_ immu_0.page_table\[4\]\[5\] _2574_ _2582_ vssd1 vssd1 vccd1 vccd1 _0148_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__5472__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7216_ clknet_leaf_22_core_clock _0477_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4428_ net89 net88 net87 net105 vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__or4b_1
XFILLER_120_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5873__A1 _2805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7147_ clknet_leaf_35_core_clock _0408_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4359_ _1523_ _1862_ _1530_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__o21a_1
XFILLER_235_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3884__A0 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7078_ clknet_leaf_11_core_clock _0339_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_219_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7399__A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6029_ _2903_ vssd1 vssd1 vccd1 vccd1 _2904_ sky130_fd_sc_hd__clkbuf_4
XFILLER_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4816__A _2166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3720__A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3964__C_N _1410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4535__B _2000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4027__S _1408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6050__A1 _2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3866__S _1386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4551__A _1910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6577__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input373_A ic1_wb_adr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input67_A c0_o_req_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6478__A _2190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5382__A _1926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4116__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6197__B _3002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5864__A1 _2618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3875__A0 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_0_0_core_clock clknet_2_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_77_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5616__A1 _2227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3627__A0 _1204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4726__A _2121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5919__A2 _2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6041__A1 _2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5395__A3 _2525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ dmmu1.page_table\[14\]\[12\] dmmu1.page_table\[15\]\[12\] _0856_ vssd1 vssd1
+ vccd1 vccd1 _1311_ sky130_fd_sc_hd__mux2_1
XANTENNA__4461__A net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3661_ dmmu0.page_table\[14\]\[11\] dmmu0.page_table\[15\]\[11\] _0896_ vssd1 vssd1
+ vccd1 vccd1 _1243_ sky130_fd_sc_hd__mux2_1
XFILLER_173_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4355__A1 _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5400_ _2310_ _2527_ vssd1 vssd1 vccd1 vccd1 _2536_ sky130_fd_sc_hd__and2_1
XFILLER_146_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6380_ net200 _3097_ vssd1 vssd1 vccd1 vccd1 _3113_ sky130_fd_sc_hd__and2_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5552__B1 _2625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3592_ dmmu0.page_table\[12\]\[9\] dmmu0.page_table\[13\]\[9\] _1169_ vssd1 vssd1
+ vccd1 vccd1 _1176_ sky130_fd_sc_hd__mux2_1
X_5331_ _2489_ immu_0.page_table\[9\]\[0\] _2495_ _2496_ vssd1 vssd1 vccd1 vccd1 _0088_
+ sky130_fd_sc_hd__a31o_1
XFILLER_142_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5292__A _2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3805__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5262_ _2447_ dmmu0.page_table\[7\]\[9\] _2445_ vssd1 vssd1 vccd1 vccd1 _2456_ sky130_fd_sc_hd__and3_1
XFILLER_272_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5855__A1 _2618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7001_ clknet_leaf_37_core_clock _0262_ vssd1 vssd1 vccd1 vccd1 immu_1.high_addr_off\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4213_ immu_0.page_table\[14\]\[7\] immu_0.page_table\[15\]\[7\] _1407_ vssd1 vssd1
+ vccd1 vccd1 _1720_ sky130_fd_sc_hd__mux2_1
XANTENNA__3866__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5193_ _2410_ vssd1 vssd1 vccd1 vccd1 _2411_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4144_ _1648_ _1651_ vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__xnor2_1
XFILLER_268_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4636__A _2054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4075_ immu_1.page_table\[14\]\[4\] immu_1.page_table\[15\]\[4\] _1438_ vssd1 vssd1
+ vccd1 vccd1 _1585_ sky130_fd_sc_hd__mux2_1
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4977_ _1987_ _2274_ _2277_ immu_1.page_table\[0\]\[9\] vssd1 vssd1 vccd1 vccd1 _0762_
+ sky130_fd_sc_hd__o22a_1
XFILLER_211_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5386__A3 _2525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5467__A _1922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4594__A1 _2019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6716_ clknet_leaf_62_core_clock _0786_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4371__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3928_ net367 vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__buf_4
XFILLER_177_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6647_ clknet_leaf_43_core_clock _0717_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3859_ net242 _1383_ net664 vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__mux2_4
XFILLER_166_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6578_ clknet_leaf_49_core_clock _0648_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4897__A2 _2219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5529_ _2603_ immu_0.page_table\[2\]\[4\] _2607_ _2613_ vssd1 vssd1 vccd1 vccd1 _0169_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__6298__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6099__A1 _2932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4310__S _1524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput560 net560 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[8] sky130_fd_sc_hd__buf_2
XFILLER_78_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5846__A1 _2618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput571 net571 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[11] sky130_fd_sc_hd__buf_2
XFILLER_160_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput582 net582 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[7] sky130_fd_sc_hd__buf_2
Xoutput593 net593 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[1] sky130_fd_sc_hd__buf_2
XFILLER_160_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5310__A3 _2480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5930__A _2834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6464__C _3159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3450__A _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6271__A1 _3042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input121_A c1_o_mem_addr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3704__S0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input219_A dcache_mem_o_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4821__A2 _2172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4034__B1 _1432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5377__A3 _2510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4585__A1 _2010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6001__A _2795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output438_A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5840__A _1968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4456__A _1940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3360__A _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4900_ _2204_ dmmu0.page_table\[0\]\[3\] _2221_ vssd1 vssd1 vccd1 vccd1 _2231_ sky130_fd_sc_hd__and3_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5880_ _2777_ dmmu0.page_table\[6\]\[0\] _2814_ vssd1 vssd1 vccd1 vccd1 _2815_ sky130_fd_sc_hd__and3_1
XFILLER_233_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4831_ net190 net189 _2027_ vssd1 vssd1 vccd1 vccd1 _2187_ sky130_fd_sc_hd__or3_2
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5287__A _2458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6892__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4762_ _2134_ immu_1.page_table\[5\]\[5\] _2140_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__and3_1
XFILLER_267_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6501_ net211 _3182_ vssd1 vssd1 vccd1 vccd1 _3183_ sky130_fd_sc_hd__or2_1
XFILLER_159_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3713_ dmmu0.page_table\[0\]\[12\] dmmu0.page_table\[1\]\[12\] net15 vssd1 vssd1
+ vccd1 vccd1 _1294_ sky130_fd_sc_hd__mux2_1
X_7481_ net178 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_2
X_4693_ _2089_ immu_1.page_table\[9\]\[0\] _2103_ vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__and3_1
X_6432_ _1898_ dmmu1.page_table\[0\]\[6\] _3135_ _3144_ vssd1 vssd1 vccd1 vccd1 _0541_
+ sky130_fd_sc_hd__a31o_1
XFILLER_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3644_ _1221_ _1226_ _0926_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__mux2_1
XANTENNA__3536__C1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6363_ net204 _3098_ vssd1 vssd1 vccd1 vccd1 _3104_ sky130_fd_sc_hd__and2_1
X_3575_ dmmu1.page_table\[0\]\[9\] dmmu1.page_table\[1\]\[9\] _0856_ vssd1 vssd1 vccd1
+ vccd1 _1159_ sky130_fd_sc_hd__mux2_1
XFILLER_136_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5540__A3 _2607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5314_ _2363_ immu_0.page_table\[10\]\[4\] _2480_ _2486_ vssd1 vssd1 vccd1 vccd1
+ _0081_ sky130_fd_sc_hd__a31o_1
XFILLER_283_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6294_ net202 _3060_ vssd1 vssd1 vccd1 vccd1 _3063_ sky130_fd_sc_hd__and2_1
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5245_ _2370_ vssd1 vssd1 vccd1 vccd1 _2447_ sky130_fd_sc_hd__clkbuf_4
XFILLER_142_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5750__A _2709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4500__A1 _1939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5176_ _2370_ vssd1 vssd1 vccd1 vccd1 _2400_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4127_ immu_0.page_table\[8\]\[6\] immu_0.page_table\[9\]\[6\] _1601_ vssd1 vssd1
+ vccd1 vccd1 _1635_ sky130_fd_sc_hd__mux2_1
XFILLER_232_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3270__A _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4058_ _1568_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4085__B immu_1.high_addr_off\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5909__B _2555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5531__A3 _2607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3445__A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6615__CLK clknet_leaf_53_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_core_clock clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_279_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input169_A c1_o_req_addr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5660__A _1896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5295__A2 _2462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input336_A ic1_mem_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6765__CLK clknet_leaf_85_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4707__C _2103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5819__B dmmu0.page_table\[3\]\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4007__B1 _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_core_clock clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_183_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output555_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3360_ _0909_ _0951_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__or2_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3291_ dmmu1.page_table\[2\]\[0\] dmmu1.page_table\[3\]\[0\] _0865_ vssd1 vssd1 vccd1
+ vccd1 _0884_ sky130_fd_sc_hd__mux2_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5286__A2 _2462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6483__A1 _1995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5030_ net103 vssd1 vssd1 vccd1 vccd1 _2310_ sky130_fd_sc_hd__buf_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6385__B _2187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3392__S1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4617__C _2049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6235__A1 _3026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6981_ clknet_leaf_78_core_clock _0242_ vssd1 vssd1 vccd1 vccd1 immu_0.high_addr_off\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_226_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7497__A net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5932_ _2834_ dmmu0.page_table\[5\]\[10\] _2831_ vssd1 vssd1 vccd1 vccd1 _2844_ sky130_fd_sc_hd__and3_1
XFILLER_280_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5863_ _2803_ _2789_ vssd1 vssd1 vccd1 vccd1 _2804_ sky130_fd_sc_hd__and2_1
XFILLER_178_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4549__A1 _2010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4814_ _2166_ immu_1.page_table\[2\]\[3\] _2174_ vssd1 vssd1 vccd1 vccd1 _2178_ sky130_fd_sc_hd__and3_1
XFILLER_33_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5794_ _2749_ dmmu0.page_table\[13\]\[8\] _2751_ vssd1 vssd1 vccd1 vccd1 _2760_ sky130_fd_sc_hd__and3_1
XFILLER_178_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5210__A2 _2409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7070__CLK clknet_leaf_4_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4745_ _2134_ immu_1.page_table\[6\]\[10\] _2122_ vssd1 vssd1 vccd1 vccd1 _2135_
+ sky130_fd_sc_hd__and3_1
XFILLER_159_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6638__CLK clknet_leaf_42_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5745__A _2731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7464_ net403 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_1
X_4676_ _2089_ immu_1.page_table\[10\]\[5\] _2086_ vssd1 vssd1 vccd1 vccd1 _2093_
+ sky130_fd_sc_hd__and3_1
XFILLER_147_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6415_ _3133_ vssd1 vssd1 vccd1 vccd1 _3134_ sky130_fd_sc_hd__clkbuf_2
XFILLER_134_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3627_ _1204_ _1209_ _0878_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__mux2_1
X_7395_ net334 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3265__A _0857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6346_ _3085_ dmmu1.page_table\[3\]\[11\] _3076_ _3092_ vssd1 vssd1 vccd1 vccd1 _0507_
+ sky130_fd_sc_hd__a31o_1
X_3558_ _1104_ _1134_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__and3_1
XANTENNA__6788__CLK clknet_leaf_2_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6277_ _3042_ dmmu1.page_table\[5\]\[9\] _3038_ _3051_ vssd1 vssd1 vccd1 vccd1 _0479_
+ sky130_fd_sc_hd__a31o_1
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3489_ _1072_ _1075_ _0899_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__mux2_1
XFILLER_276_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5480__A net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput107 c1_o_c_instr_long vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_4
Xinput118 c1_o_mem_addr[0] vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__buf_2
X_5228_ _1913_ _2350_ vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__nor2_2
XANTENNA__5911__C _2832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput129 c1_o_mem_addr[5] vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_2
XFILLER_229_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5159_ _2389_ vssd1 vssd1 vccd1 vccd1 _2390_ sky130_fd_sc_hd__buf_4
XANTENNA__3383__S1 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6226__A1 _3010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_2_1_0_core_clock_A clknet_1_0_1_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3460__A1 _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5201__A2 _2409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input286_A ic0_mem_data[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5374__B _2512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5504__A3 _2591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4712__A1 _2021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6465__A1 _1974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3374__S1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_57_core_clock_A clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__6217__A1 _3010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4734__A _2121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7093__CLK clknet_leaf_32_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3451__A1 _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output672_A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4400__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4530_ _1995_ vssd1 vssd1 vccd1 vccd1 _1996_ sky130_fd_sc_hd__buf_6
XANTENNA__4951__A1 _1979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4900__C _2221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4461_ net102 vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__buf_4
XFILLER_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6200_ _2994_ dmmu1.page_table\[7\]\[3\] _3000_ _3006_ vssd1 vssd1 vccd1 vccd1 _0447_
+ sky130_fd_sc_hd__a31o_1
X_3412_ dmmu1.page_table\[0\]\[4\] dmmu1.page_table\[1\]\[4\] dmmu1.page_table\[2\]\[4\]
+ dmmu1.page_table\[3\]\[4\] _0865_ _0863_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__mux4_1
XANTENNA__4164__C1 _1553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7180_ clknet_leaf_29_core_clock _0441_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[8\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4392_ net272 _1892_ _0811_ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__mux2_4
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _2845_ dmmu0.page_table\[1\]\[2\] _2962_ vssd1 vssd1 vccd1 vccd1 _2965_ sky130_fd_sc_hd__and3_1
X_3343_ dmmu1.page_table\[8\]\[1\] dmmu1.page_table\[9\]\[1\] dmmu1.page_table\[10\]\[1\]
+ dmmu1.page_table\[11\]\[1\] _0891_ _0860_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__mux4_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4909__A _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5259__A2 _2442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6062_ _2923_ vssd1 vssd1 vccd1 vccd1 _2924_ sky130_fd_sc_hd__clkbuf_4
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3274_ _0864_ _0866_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__or2_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _1897_ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__buf_4
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6964_ clknet_leaf_90_core_clock _0225_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5459__B _2559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5915_ _2223_ _2830_ _2835_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__a21o_1
X_6895_ clknet_leaf_71_core_clock _0156_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5846_ _2618_ dmmu1.page_table\[15\]\[1\] _2787_ _2792_ vssd1 vssd1 vccd1 vccd1 _0307_
+ sky130_fd_sc_hd__a31o_1
XFILLER_42_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5195__A1 _2211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5777_ _2750_ vssd1 vssd1 vccd1 vccd1 _2751_ sky130_fd_sc_hd__buf_2
XFILLER_194_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4942__A1 _1967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4728_ _2121_ immu_1.page_table\[6\]\[2\] _2123_ vssd1 vssd1 vccd1 vccd1 _2126_ sky130_fd_sc_hd__and3_1
XFILLER_135_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4810__C _2174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7447_ net61 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_1
X_4659_ _1959_ _2062_ vssd1 vssd1 vccd1 vccd1 _2081_ sky130_fd_sc_hd__or2_4
XFILLER_206_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7378_ net710 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_1
XFILLER_89_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6329_ _3069_ dmmu1.page_table\[3\]\[3\] _3077_ _3083_ vssd1 vssd1 vccd1 vccd1 _0499_
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6447__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_5_0_core_clock clknet_2_2_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3681__A1 _0868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3869__S _1390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4554__A _1910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6803__CLK clknet_leaf_81_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6472__C _3159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input201_A c1_sr_bus_data_o[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5973__A3 _2859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5186__A1 _2251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input97_A c0_sr_bus_data_o[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5385__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4933__A1 _2253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7309__CLK clknet_leaf_19_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5832__B dmmu0.page_table\[3\]\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6438__A1 _1898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output518_A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3672__B2 _0957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4464__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3961_ immu_0.page_table\[2\]\[1\] immu_0.page_table\[3\]\[1\] _1407_ vssd1 vssd1
+ vccd1 vccd1 _1474_ sky130_fd_sc_hd__mux2_1
XANTENNA__5964__A3 _2859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5700_ _2682_ dmmu0.page_table\[2\]\[3\] _2702_ vssd1 vssd1 vccd1 vccd1 _2706_ sky130_fd_sc_hd__and3_1
XFILLER_259_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6680_ clknet_leaf_54_core_clock _0750_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[7\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3892_ _1406_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_1
XFILLER_189_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5631_ _2655_ dmmu0.page_table\[15\]\[10\] _2651_ vssd1 vssd1 vccd1 vccd1 _2664_
+ sky130_fd_sc_hd__and3_1
X_5562_ _2628_ vssd1 vssd1 vccd1 vccd1 _2629_ sky130_fd_sc_hd__inv_2
XANTENNA__4924__A1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7301_ clknet_leaf_44_core_clock _0562_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[8\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4513_ _1976_ dmmu1.page_table\[14\]\[7\] _1964_ _1984_ vssd1 vssd1 vccd1 vccd1 _0591_
+ sky130_fd_sc_hd__a31o_1
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5493_ _2588_ immu_0.page_table\[3\]\[0\] _2591_ _2592_ vssd1 vssd1 vccd1 vccd1 _0154_
+ sky130_fd_sc_hd__a31o_1
X_7232_ clknet_leaf_27_core_clock _0493_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[4\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4444_ _1911_ immu_0.page_table\[11\]\[1\] _1924_ _1932_ vssd1 vssd1 vccd1 vccd1
+ _0574_ sky130_fd_sc_hd__a31o_1
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5742__B _2572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7163_ clknet_leaf_9_core_clock _0424_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4375_ net107 _1877_ _1878_ vssd1 vssd1 vccd1 vccd1 _1879_ sky130_fd_sc_hd__and3_1
X_6114_ _2948_ dmmu1.page_table\[9\]\[8\] _2942_ _2954_ vssd1 vssd1 vccd1 vccd1 _0413_
+ sky130_fd_sc_hd__a31o_1
X_3326_ dmmu0.page_table\[8\]\[0\] dmmu0.page_table\[9\]\[0\] dmmu0.page_table\[10\]\[0\]
+ dmmu0.page_table\[11\]\[0\] _0897_ _0902_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__mux4_1
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7094_ clknet_leaf_11_core_clock _0355_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_219_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6045_ _2898_ dmmu1.page_table\[11\]\[7\] _2902_ _2912_ vssd1 vssd1 vccd1 vccd1 _0386_
+ sky130_fd_sc_hd__a31o_1
XFILLER_218_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3257_ net133 net28 _0847_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__mux2_2
XFILLER_273_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3188_ _0811_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_12
XANTENNA__3689__S _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3415__A1 _0881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6947_ clknet_leaf_1_core_clock _0208_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[12\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_241_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3510__S1 _0902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6878_ clknet_leaf_71_core_clock _0139_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5829_ _1948_ _2767_ _2780_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__a21o_1
XFILLER_167_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4376__C1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5340__A1 _2489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3453__A _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input151_A c1_o_mem_high_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input249_A dcache_wb_adr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5643__A2 _2669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4300__C1 _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3599__S _1169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input12_A c0_o_instr_long_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4284__A _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output468_A net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5331__A1 _2489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output635_A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4459__A _1942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4160_ immu_1.page_table\[0\]\[6\] immu_1.page_table\[1\]\[6\] _1438_ vssd1 vssd1
+ vccd1 vccd1 _1668_ sky130_fd_sc_hd__mux2_1
XANTENNA__5281__C _2464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4091_ immu_0.page_table\[4\]\[5\] immu_0.page_table\[5\]\[5\] immu_0.page_table\[6\]\[5\]
+ immu_0.page_table\[7\]\[5\] _1409_ _1570_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__mux4_2
XFILLER_67_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6999__CLK clknet_leaf_38_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput290 ic0_mem_data[21] vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_1
XANTENNA__6393__B _3118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3645__B2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4842__B1 _2192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4625__C _2049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6801_ clknet_leaf_6_core_clock _0062_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[7\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4993_ _2284_ immu_1.page_table\[15\]\[4\] _2282_ vssd1 vssd1 vccd1 vccd1 _2288_
+ sky130_fd_sc_hd__and3_1
XFILLER_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6732_ clknet_leaf_63_core_clock _0802_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4922__A _1948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3944_ _1445_ _1452_ _1455_ _1456_ _1457_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__o221a_1
XANTENNA__4070__A1 _1411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6663_ clknet_leaf_9_core_clock _0733_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3875_ net321 net375 _1390_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__mux2_1
XFILLER_149_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3538__A net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5614_ _2370_ vssd1 vssd1 vccd1 vccd1 _2655_ sky130_fd_sc_hd__clkbuf_4
XFILLER_136_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6594_ clknet_leaf_54_core_clock _0664_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_219_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6362__A3 _3096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5545_ _2622_ vssd1 vssd1 vccd1 vccd1 _2623_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5570__A1 _2239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3972__S _1443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5753__A _2736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5476_ net100 _2577_ vssd1 vssd1 vccd1 vccd1 _2582_ sky130_fd_sc_hd__and2_1
XFILLER_144_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6114__A3 _2942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5472__B _2577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7215_ clknet_leaf_14_core_clock _0476_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4427_ _1915_ _1916_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__or2_1
XFILLER_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7146_ clknet_leaf_14_core_clock _0407_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4358_ immu_1.page_table\[10\]\[10\] immu_1.page_table\[11\]\[10\] _1439_ vssd1 vssd1
+ vccd1 vccd1 _1862_ sky130_fd_sc_hd__mux2_1
XANTENNA__3884__A1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input4_A c0_o_icache_flush vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3309_ _0901_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__buf_4
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7077_ clknet_leaf_78_core_clock _0338_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4289_ _1570_ _1791_ _1793_ _1535_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__o211a_1
XFILLER_274_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6028_ _1968_ _2064_ vssd1 vssd1 vccd1 vccd1 _2903_ sky130_fd_sc_hd__nor2_1
XFILLER_104_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7004__CLK clknet_leaf_36_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7154__CLK clknet_leaf_29_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5928__A _2834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4832__A _1999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3495__S0 _0858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input199_A c1_sr_bus_data_o[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3882__S _1386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input366_A ic1_wb_adr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3875__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3911__A _1407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5616__A2 _2650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4218__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5092__A3 _2336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4742__A _2121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4052__A1 _1523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3486__S0 _0900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6521__CLK clknet_leaf_43_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3660_ _0909_ _1239_ _1241_ _0917_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__o211a_1
XFILLER_9_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5552__A1 _2232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3591_ _0912_ _1174_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__nand2_1
XANTENNA__6671__CLK clknet_leaf_4_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5330_ _1926_ _2494_ vssd1 vssd1 vccd1 vccd1 _2496_ sky130_fd_sc_hd__nor2_1
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3805__B _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5261_ _2245_ _2442_ _2455_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__a21o_1
XFILLER_114_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7000_ clknet_leaf_37_core_clock _0261_ vssd1 vssd1 vccd1 vccd1 immu_1.high_addr_off\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4212_ _1430_ _1716_ _1718_ _1416_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__o211a_1
XFILLER_141_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5192_ _2216_ _2407_ vssd1 vssd1 vccd1 vccd1 _2410_ sky130_fd_sc_hd__or2_1
XANTENNA__3410__S0 _0891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3866__A1 _1388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4143_ _1649_ _1650_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__and2b_1
XFILLER_228_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4917__A _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3821__A inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4074_ _1446_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__buf_2
XFILLER_83_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7177__CLK clknet_leaf_33_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5083__A3 _2336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5748__A _2709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4976_ _1985_ _2274_ _2277_ immu_1.page_table\[0\]\[8\] vssd1 vssd1 vccd1 vccd1 _0761_
+ sky130_fd_sc_hd__o22a_1
XFILLER_51_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5467__B _2572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6715_ clknet_leaf_61_core_clock _0785_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[15\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4594__A2 _2030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5791__A1 _2239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3927_ net385 net108 _1440_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__and3b_2
XANTENNA__3268__A _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6646_ clknet_leaf_42_core_clock _0716_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3858_ net316 net370 _1360_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__mux2_2
XFILLER_177_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6577_ clknet_leaf_49_core_clock _0647_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3789_ _1345_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_31_core_clock clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5914__C _2832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5528_ net99 _2609_ vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__and2_1
XANTENNA__6298__B _3060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5459_ _2314_ _2559_ vssd1 vssd1 vccd1 vccd1 _2571_ sky130_fd_sc_hd__and2_1
Xoutput550 net550 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[13] sky130_fd_sc_hd__buf_2
Xoutput561 net561 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[9] sky130_fd_sc_hd__buf_2
XFILLER_105_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput572 net572 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[12] sky130_fd_sc_hd__buf_2
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput583 net583 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[8] sky130_fd_sc_hd__buf_2
XFILLER_266_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput594 net594 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[2] sky130_fd_sc_hd__buf_2
XFILLER_59_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7129_ clknet_leaf_29_core_clock _0390_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[11\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_219_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4827__A _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3609__A1 _0929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3609__B2 _0957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3704__S1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6544__CLK clknet_leaf_50_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input114_A c1_o_instr_long_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5658__A _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4034__A1 _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5231__B1 _1911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4585__A2 _2030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_core_clock clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_230_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6694__CLK clknet_leaf_41_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3906__A _1419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6001__B _2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5840__B _2278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4456__B _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4273__A1 _1516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4830_ _2025_ _2171_ _2186_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__a21o_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4761_ _2012_ _2138_ _2145_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__a21o_1
XFILLER_221_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3712_ dmmu0.page_table\[2\]\[12\] dmmu0.page_table\[3\]\[12\] net15 vssd1 vssd1
+ vccd1 vccd1 _1293_ sky130_fd_sc_hd__mux2_1
X_6500_ net96 icore_sregs.c1_disable _3181_ vssd1 vssd1 vccd1 vccd1 _3182_ sky130_fd_sc_hd__mux2_1
XFILLER_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7480_ net177 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__buf_2
XFILLER_159_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4692_ _2102_ vssd1 vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__buf_2
XFILLER_201_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6431_ net206 _3137_ vssd1 vssd1 vccd1 vccd1 _3144_ sky130_fd_sc_hd__and2_1
XANTENNA__5525__A1 _2603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3643_ _1224_ _1225_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__xnor2_1
XANTENNA__6399__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6362_ _3101_ dmmu1.page_table\[2\]\[3\] _3096_ _3103_ vssd1 vssd1 vccd1 vccd1 _0512_
+ sky130_fd_sc_hd__a31o_1
XFILLER_283_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3574_ dmmu1.page_table\[2\]\[9\] dmmu1.page_table\[3\]\[9\] _0857_ vssd1 vssd1 vccd1
+ vccd1 _1158_ sky130_fd_sc_hd__mux2_1
XFILLER_127_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5313_ _1937_ _2482_ vssd1 vssd1 vccd1 vccd1 _2486_ sky130_fd_sc_hd__and2_1
XFILLER_161_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6293_ _3053_ dmmu1.page_table\[4\]\[1\] _3058_ _3062_ vssd1 vssd1 vccd1 vccd1 _0484_
+ sky130_fd_sc_hd__a31o_1
XFILLER_102_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5244_ _2211_ _2442_ _2446_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__a21o_1
XFILLER_142_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4647__A _2072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5175_ _2240_ _2390_ _2399_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__a21o_1
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4126_ _1569_ net239 _1614_ _1634_ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__a22o_4
XFILLER_256_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6567__CLK clknet_leaf_50_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5056__A3 _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4057_ net237 _1567_ _0811_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__mux2_1
XFILLER_271_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5478__A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4382__A _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4016__A1 _1523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5764__A1 _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4959_ _1987_ _2257_ _2270_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__a21o_1
XFILLER_177_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6308__A3 _3058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6629_ clknet_leaf_56_core_clock _0699_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_257_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6102__A _2931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5644__C _2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4557__A _1897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input231_A dcache_wb_adr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input329_A ic0_wb_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4007__A1 _1448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3766__A0 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4231__S _1601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6012__A _2891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6180__A1 _2977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3613__S0 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output450_A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output548_A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5851__A _2795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3290_ _0864_ _0882_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__or2_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4467__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4494__A1 _1939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6980_ clknet_leaf_78_core_clock _0241_ vssd1 vssd1 vccd1 vccd1 immu_0.high_addr_off\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_253_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5931_ _1948_ _2830_ _2843_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__a21o_1
XFILLER_213_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5298__A _2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5862_ net207 vssd1 vssd1 vccd1 vccd1 _2803_ sky130_fd_sc_hd__clkbuf_4
XFILLER_278_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4549__A2 _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4813_ _2008_ _2172_ _2177_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__a21o_1
X_5793_ _2242_ _2748_ _2759_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__a21o_1
XFILLER_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4744_ _2105_ vssd1 vssd1 vccd1 vccd1 _2134_ sky130_fd_sc_hd__clkbuf_4
XFILLER_119_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4675_ _2012_ _2083_ _2092_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__a21o_1
X_7463_ net402 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_1
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3509__B1 _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6414_ _1958_ _2272_ vssd1 vssd1 vccd1 vccd1 _3133_ sky130_fd_sc_hd__or2_1
X_3626_ _1207_ _1208_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__xor2_1
X_7394_ net333 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_1
XFILLER_162_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6345_ net199 _3078_ vssd1 vssd1 vccd1 vccd1 _3092_ sky130_fd_sc_hd__and2_1
X_3557_ _0921_ _1137_ _1141_ _0957_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__a211o_1
XANTENNA__5761__A _2736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6276_ _2893_ _3040_ vssd1 vssd1 vccd1 vccd1 _3051_ sky130_fd_sc_hd__and2_1
X_3488_ _1073_ _1074_ _0917_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__mux2_1
XFILLER_88_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5480__B _2577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5227_ _2210_ _2428_ _2431_ vssd1 vssd1 vccd1 vccd1 _2432_ sky130_fd_sc_hd__a21oi_1
Xinput108 c1_o_c_instr_page vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_2
Xinput119 c1_o_mem_addr[10] vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__buf_2
XFILLER_130_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4377__A inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3281__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5682__A0 _2232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4808__C _2174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5158_ _2217_ _2388_ vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__nor2_1
XFILLER_56_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5029__A3 _2298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4109_ _1615_ _1616_ _1596_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__a21boi_1
XFILLER_229_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5089_ _2332_ immu_0.page_table\[12\]\[8\] _2336_ _2346_ vssd1 vssd1 vccd1 vccd1
+ _0805_ sky130_fd_sc_hd__a31o_1
XFILLER_217_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5985__A1 _2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3996__B1 _1479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5001__A _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4096__S0 _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3748__A0 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input181_A c1_sr_bus_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6162__A1 _2977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input279_A ic0_mem_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6732__CLK clknet_leaf_63_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4173__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4712__A2 _2101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3890__S _1390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5671__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input42_A c0_o_mem_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6465__A2 _3157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6882__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3191__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5440__A3 _2557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6007__A _2801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5728__A1 _1967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3739__A0 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4750__A _2084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4400__A1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4951__A2 _2257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3366__A _0957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4460_ _1939_ immu_0.page_table\[11\]\[6\] _1924_ _1943_ vssd1 vssd1 vccd1 vccd1
+ _0579_ sky130_fd_sc_hd__a31o_1
XANTENNA__6153__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3411_ _0855_ _0999_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__or2_1
XFILLER_144_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5900__A1 _1948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4391_ net326 net380 _0812_ vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__mux2_2
XFILLER_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5581__A _2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6130_ _2223_ _2960_ _2964_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__a21o_1
X_3342_ _0869_ _0931_ _0933_ _0854_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__o211a_1
XFILLER_98_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__B _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6061_ _1968_ _2081_ vssd1 vssd1 vccd1 vccd1 _2923_ sky130_fd_sc_hd__nor2_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4197__A _1457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3273_ dmmu1.page_table\[8\]\[0\] dmmu1.page_table\[9\]\[0\] _0865_ vssd1 vssd1 vccd1
+ vccd1 _0866_ sky130_fd_sc_hd__mux2_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5012_ _1976_ immu_0.page_table\[15\]\[0\] _2298_ _2299_ vssd1 vssd1 vccd1 vccd1
+ _0775_ sky130_fd_sc_hd__a31o_1
XFILLER_285_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4925__A _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6963_ clknet_leaf_88_core_clock _0224_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_241_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5914_ _2834_ dmmu0.page_table\[5\]\[1\] _2832_ vssd1 vssd1 vccd1 vccd1 _2835_ sky130_fd_sc_hd__and3_1
XANTENNA__6605__CLK clknet_leaf_54_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6894_ clknet_leaf_72_core_clock _0155_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5845_ _2791_ _2789_ vssd1 vssd1 vccd1 vccd1 _2792_ sky130_fd_sc_hd__and2_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4660__A _2000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5195__A2 _2409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6392__A1 _3112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5776_ _2443_ _2351_ vssd1 vssd1 vccd1 vccd1 _2750_ sky130_fd_sc_hd__or2_2
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4727_ _2006_ _2120_ _2125_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__a21o_1
XANTENNA__4942__A2 _2257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3276__A _0868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5194__C _2411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7446_ net60 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_1
XFILLER_174_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4658_ _2025_ _2065_ _2080_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__a21o_1
XFILLER_162_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput90 c0_sr_bus_addr[8] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5498__A3 _2591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3609_ _0929_ _1178_ _1187_ _1192_ _0957_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__a32o_1
X_7377_ net276 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_2
X_4589_ _2038_ immu_1.page_table\[13\]\[5\] _2032_ vssd1 vssd1 vccd1 vccd1 _2039_
+ sky130_fd_sc_hd__and3_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5922__C _2832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6328_ net203 _3079_ vssd1 vssd1 vccd1 vccd1 _3083_ sky130_fd_sc_hd__and2_1
XFILLER_107_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6447__A2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6259_ _2931_ vssd1 vssd1 vccd1 vccd1 _3042_ sky130_fd_sc_hd__buf_4
XFILLER_276_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4835__A _2190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5422__A3 _2541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3969__B1 _1411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4046__S _1443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3885__S _1386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5666__A _2682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4570__A _2017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input396_A inner_wb_i_dat[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4394__A0 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5385__B _2527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4146__B1 _1653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7060__CLK clknet_leaf_79_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4745__A _2134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5413__A3 _2541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5279__C _2464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3960_ immu_0.page_table\[4\]\[1\] immu_0.page_table\[5\]\[1\] immu_0.page_table\[6\]\[1\]
+ immu_0.page_table\[7\]\[1\] _1472_ _1419_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__mux4_2
XANTENNA__6778__CLK clknet_leaf_85_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3891_ net233 _1405_ _1386_ vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__mux2_4
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3975__A3 immu_1.page_table\[7\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4480__A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5630_ _2247_ _2650_ _2663_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__a21o_1
XFILLER_176_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6374__A1 _3101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4385__B1 _1360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5561_ _2190_ _2626_ vssd1 vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__nand2_1
XANTENNA__4924__A2 _2219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7300_ clknet_leaf_44_core_clock _0561_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[8\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4512_ _1983_ _1970_ vssd1 vssd1 vccd1 vccd1 _1984_ sky130_fd_sc_hd__and2_1
X_5492_ _1925_ _2590_ vssd1 vssd1 vccd1 vccd1 _2592_ sky130_fd_sc_hd__nor2_1
XFILLER_156_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7231_ clknet_leaf_23_core_clock _0492_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[4\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_4443_ _1928_ _1931_ vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__and2_1
XFILLER_208_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3824__A _1363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7162_ clknet_leaf_11_core_clock _0423_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4374_ _1806_ _1876_ _1875_ _1874_ vssd1 vssd1 vccd1 vccd1 _1878_ sky130_fd_sc_hd__o211ai_1
XFILLER_258_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6113_ _2891_ _2944_ vssd1 vssd1 vccd1 vccd1 _2954_ sky130_fd_sc_hd__and2_1
X_3325_ _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__buf_4
X_7093_ clknet_leaf_32_core_clock _0354_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6044_ _2803_ _2904_ vssd1 vssd1 vccd1 vccd1 _2912_ sky130_fd_sc_hd__and2_1
X_3256_ _0851_ vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4655__A _2072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3187_ inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__inv_6
XFILLER_226_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4860__A1 _1974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6946_ clknet_leaf_81_core_clock _0207_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[12\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_240_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6877_ clknet_leaf_70_core_clock _0138_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5486__A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4390__A _1891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5828_ _2777_ dmmu0.page_table\[3\]\[9\] _2769_ vssd1 vssd1 vccd1 vccd1 _2780_ sky130_fd_sc_hd__and3_1
XFILLER_167_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5759_ _2736_ dmmu0.page_table\[4\]\[6\] _2732_ vssd1 vssd1 vccd1 vccd1 _2740_ sky130_fd_sc_hd__and3_1
XFILLER_108_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7429_ net390 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_1
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4679__A1 _2016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5652__C _2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7083__CLK clknet_leaf_5_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input144_A c1_o_mem_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4300__B1 _1804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input311_A ic0_wb_adr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6920__CLK clknet_leaf_76_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5396__A _1942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3909__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6108__A1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_69_core_clock_A clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_99_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6020__A _1991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4459__B _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3342__A1 _0869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output530_A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output628_A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4090_ _1569_ net238 _1580_ _1599_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__a22o_4
XFILLER_255_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput280 ic0_mem_data[12] vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4842__A1 _1979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput291 ic0_mem_data[22] vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_1
XFILLER_208_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6800_ clknet_leaf_6_core_clock _0061_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[7\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4992_ _1974_ _2280_ _2287_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__a21o_1
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6731_ clknet_leaf_67_core_clock _0801_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_223_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3943_ net369 vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__clkinv_4
XFILLER_210_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4070__A2 _1575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6662_ clknet_leaf_80_core_clock _0732_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3874_ _1394_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__clkbuf_1
X_5613_ _2224_ _2650_ _2654_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__a21o_1
X_6593_ clknet_leaf_59_core_clock _0663_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_117_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5544_ _1921_ _2621_ vssd1 vssd1 vccd1 vccd1 _2622_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_21_core_clock clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5475_ _2576_ immu_0.page_table\[4\]\[4\] _2574_ _2581_ vssd1 vssd1 vccd1 vccd1 _0147_
+ sky130_fd_sc_hd__a31o_1
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7214_ clknet_leaf_15_core_clock _0475_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4426_ net78 net77 net91 net90 vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__or4b_1
XFILLER_259_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7145_ clknet_leaf_33_core_clock _0406_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4357_ _1496_ _1860_ vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__or2_1
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3308_ net16 vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__clkbuf_4
XFILLER_86_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4288_ _1424_ _1792_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__or2_1
X_7076_ clknet_leaf_79_core_clock _0337_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6943__CLK clknet_leaf_85_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6027_ _2901_ vssd1 vssd1 vccd1 vccd1 _2902_ sky130_fd_sc_hd__buf_4
X_3239_ _0842_ vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_71_core_clock_A clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4816__C _2174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6050__A3 _2902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6929_ clknet_leaf_77_core_clock _0190_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4832__B _2187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3495__S1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_core_clock clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__6105__A _2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6338__A1 _3085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4551__C _2004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input261_A dcache_wb_o_dat[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input359_A ic1_mem_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5864__A3 _2787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5077__A1 _2332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4824__A1 _2019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4285__C1 _1479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4726__C _2123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6041__A3 _2902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3486__S1 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6329__A1 _3069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6015__A _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5854__A _2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3590_ dmmu0.page_table\[14\]\[9\] dmmu0.page_table\[15\]\[9\] _1169_ vssd1 vssd1
+ vccd1 vccd1 _1174_ sky130_fd_sc_hd__mux2_1
XANTENNA__5552__A2 _2623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5292__C _2464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5260_ _2447_ dmmu0.page_table\[7\]\[8\] _2445_ vssd1 vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__and3_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6966__CLK clknet_leaf_86_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4211_ _1423_ _1717_ vssd1 vssd1 vccd1 vccd1 _1718_ sky130_fd_sc_hd__or2_1
XFILLER_102_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5855__A3 _2787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5191_ _2408_ vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__buf_4
XFILLER_68_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3410__S1 _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4142_ net7 immu_0.high_addr_off\[2\] vssd1 vssd1 vccd1 vccd1 _1650_ sky130_fd_sc_hd__nand2_1
XFILLER_256_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4073_ immu_1.page_table\[12\]\[4\] immu_1.page_table\[13\]\[4\] _1439_ vssd1 vssd1
+ vccd1 vccd1 _1583_ sky130_fd_sc_hd__mux2_1
XFILLER_228_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4815__A1 _2010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4636__C _2068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4975_ _1983_ _2274_ _2277_ immu_1.page_table\[0\]\[7\] vssd1 vssd1 vccd1 vccd1 _0760_
+ sky130_fd_sc_hd__o22a_1
XFILLER_211_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3251__A0 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6714_ clknet_leaf_62_core_clock _0784_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[15\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3926_ net107 vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__clkinv_2
XFILLER_211_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5791__A2 _2748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6645_ clknet_leaf_40_core_clock _0715_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3857_ _1382_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6576_ clknet_leaf_46_core_clock _0646_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3788_ net223 _0993_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__and2_1
XFILLER_119_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5527_ _2603_ immu_0.page_table\[2\]\[3\] _2607_ _2612_ vssd1 vssd1 vccd1 vccd1 _0168_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__3284__A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6099__A3 _2942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5458_ _2562_ immu_0.page_table\[5\]\[9\] _2557_ _2570_ vssd1 vssd1 vccd1 vccd1 _0141_
+ sky130_fd_sc_hd__a31o_1
Xoutput540 net540 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[5] sky130_fd_sc_hd__buf_2
XFILLER_172_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput551 net551 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[14] sky130_fd_sc_hd__buf_2
Xoutput562 net562 vssd1 vssd1 vccd1 vccd1 dcache_mem_req sky130_fd_sc_hd__buf_2
XFILLER_278_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5846__A3 _2787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput573 net573 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[13] sky130_fd_sc_hd__buf_2
XFILLER_120_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4409_ _1904_ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_1
Xoutput584 net584 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[9] sky130_fd_sc_hd__buf_2
XFILLER_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput595 net595 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[3] sky130_fd_sc_hd__buf_2
X_5389_ _1935_ _2527_ vssd1 vssd1 vccd1 vccd1 _2530_ sky130_fd_sc_hd__and2_1
XFILLER_132_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7128_ clknet_leaf_29_core_clock _0389_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[11\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5930__C _2832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7059_ clknet_leaf_80_core_clock _0320_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__7121__CLK clknet_leaf_13_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3609__A2 _1178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6271__A3 _3038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4019__C1 _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7271__CLK clknet_leaf_25_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input107_A c1_o_c_instr_long vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3459__A _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6839__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3242__A0 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input72_A c0_o_req_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6989__CLK clknet_leaf_7_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5287__C _2464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _2134_ immu_1.page_table\[5\]\[4\] _2140_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__and3_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3711_ dmmu0.page_table\[4\]\[12\] dmmu0.page_table\[5\]\[12\] dmmu0.page_table\[6\]\[12\]
+ dmmu0.page_table\[7\]\[12\] _0895_ net16 vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__mux4_1
XFILLER_267_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4691_ _2084_ _2099_ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__or2_1
XFILLER_159_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6430_ _3128_ dmmu1.page_table\[0\]\[5\] _3135_ _3143_ vssd1 vssd1 vccd1 vccd1 _0540_
+ sky130_fd_sc_hd__a31o_1
X_3642_ _1189_ _1191_ _1188_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__a21bo_1
XFILLER_174_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6399__B _3118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3536__B2 _0881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6361_ net203 _3098_ vssd1 vssd1 vccd1 vccd1 _3103_ sky130_fd_sc_hd__and2_1
X_3573_ _0859_ _1156_ _0872_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__a21o_1
XFILLER_283_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5312_ _2363_ immu_0.page_table\[10\]\[3\] _2480_ _2485_ vssd1 vssd1 vccd1 vccd1
+ _0080_ sky130_fd_sc_hd__a31o_1
X_6292_ net201 _3060_ vssd1 vssd1 vccd1 vccd1 _3062_ sky130_fd_sc_hd__and2_1
XFILLER_88_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5243_ _2416_ dmmu0.page_table\[7\]\[0\] _2445_ vssd1 vssd1 vccd1 vccd1 _2446_ sky130_fd_sc_hd__and3_1
XFILLER_216_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7144__CLK clknet_leaf_34_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4928__A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3832__A _1363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3395__S0 _0898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5750__C _2732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5174_ _2384_ dmmu0.page_table\[9\]\[6\] _2392_ vssd1 vssd1 vccd1 vccd1 _2399_ sky130_fd_sc_hd__and3_1
XANTENNA__4500__A3 _1964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4125_ _1569_ _1633_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__nor2_1
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4249__C1 _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7294__CLK clknet_leaf_43_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4056_ _1552_ _1566_ _1390_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__mux2_1
XFILLER_209_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5759__A _2736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4663__A _2084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5478__B _2577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4958_ _2262_ immu_1.page_table\[7\]\[9\] _2259_ vssd1 vssd1 vccd1 vccd1 _2270_ sky130_fd_sc_hd__and3_1
XANTENNA__5764__A2 _2730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3909_ net313 vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__clkinv_2
XANTENNA__4972__B1 _2277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4889_ _2211_ _2219_ _2222_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__a21o_1
XANTENNA__5494__A _1922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6628_ clknet_leaf_55_core_clock _0698_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_257_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3527__A1 _1087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6559_ clknet_leaf_48_core_clock _0629_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[12\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_152_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3742__A _1320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6511__CLK clknet_leaf_59_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4049__S _1493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input224_A dcache_mem_o_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5452__A1 _2562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3888__S _1386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6661__CLK clknet_leaf_80_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__A1 _2233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3310__S0 _0900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6012__B _2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7167__CLK clknet_leaf_4_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3613__S1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5851__B _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output443_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4748__A _2000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3377__S0 _0898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6235__A3 _3019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5579__A _2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4483__A _1958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5930_ _2834_ dmmu0.page_table\[5\]\[9\] _2832_ vssd1 vssd1 vccd1 vccd1 _2843_ sky130_fd_sc_hd__and3_1
XFILLER_206_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5861_ _2618_ dmmu1.page_table\[15\]\[6\] _2787_ _2802_ vssd1 vssd1 vccd1 vccd1 _0312_
+ sky130_fd_sc_hd__a31o_1
XFILLER_202_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4812_ _2166_ immu_1.page_table\[2\]\[2\] _2174_ vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__and3_1
X_5792_ _2749_ dmmu0.page_table\[13\]\[7\] _2751_ vssd1 vssd1 vccd1 vccd1 _2759_ sky130_fd_sc_hd__and3_1
XFILLER_178_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4743_ _2023_ _2120_ _2133_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__a21o_1
XFILLER_193_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7462_ net401 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__clkbuf_1
XANTENNA__6203__A _2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4674_ _2089_ immu_1.page_table\[10\]\[4\] _2086_ vssd1 vssd1 vccd1 vccd1 _2092_
+ sky130_fd_sc_hd__and3_1
X_6413_ _3128_ dmmu1.page_table\[1\]\[12\] _3115_ _3132_ vssd1 vssd1 vccd1 vccd1 _0534_
+ sky130_fd_sc_hd__a31o_1
X_3625_ _1164_ _1166_ _1163_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__a21boi_1
X_7393_ net332 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_1
XFILLER_227_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6344_ _3085_ dmmu1.page_table\[3\]\[10\] _3076_ _3091_ vssd1 vssd1 vccd1 vccd1 _0506_
+ sky130_fd_sc_hd__a31o_1
X_3556_ _0899_ _1140_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__and2_1
XFILLER_115_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6275_ _3042_ dmmu1.page_table\[5\]\[8\] _3038_ _3050_ vssd1 vssd1 vccd1 vccd1 _0478_
+ sky130_fd_sc_hd__a31o_1
X_3487_ dmmu0.page_table\[8\]\[6\] dmmu0.page_table\[9\]\[6\] dmmu0.page_table\[10\]\[6\]
+ dmmu0.page_table\[11\]\[6\] _0900_ _0912_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__mux4_1
XFILLER_170_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3562__A _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5226_ net197 _2430_ net407 vssd1 vssd1 vccd1 vccd1 _2431_ sky130_fd_sc_hd__a21bo_1
Xinput109 c1_o_icache_flush vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_2
XFILLER_276_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4377__B net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_core_clock_A clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6684__CLK clknet_leaf_42_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5157_ _1913_ _2350_ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__or2_4
XFILLER_84_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4108_ _1596_ _1615_ _1616_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__and3b_1
XANTENNA__6226__A3 _3019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5088_ _2310_ _2338_ vssd1 vssd1 vccd1 vccd1 _2346_ sky130_fd_sc_hd__and2_1
XFILLER_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4393__A _1893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4039_ _1423_ _1547_ _1549_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__a21o_1
XFILLER_232_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3996__A1 _1411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4096__S1 _1570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4332__S _1480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6113__A _2891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4173__A1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input174_A c1_o_req_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input341_A ic1_mem_data[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3191__B _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_A c0_o_mem_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4734__C _2123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6007__B _2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4750__B _2136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3647__A _1229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6023__A _1993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6557__CLK clknet_leaf_48_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output560_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3410_ dmmu1.page_table\[8\]\[4\] dmmu1.page_table\[9\]\[4\] dmmu1.page_table\[10\]\[4\]
+ dmmu1.page_table\[11\]\[4\] _0891_ _0860_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__mux4_1
XANTENNA__4164__A1 _1516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4390_ _1891_ vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_1
XFILLER_264_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5900__A2 _2812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3341_ _0863_ _0932_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__or2_1
XANTENNA__4478__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4909__C _2221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _2921_ vssd1 vssd1 vccd1 vccd1 _2922_ sky130_fd_sc_hd__buf_4
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3272_ _0857_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__buf_6
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_1_core_clock_A clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _1926_ _2297_ vssd1 vssd1 vccd1 vccd1 _2299_ sky130_fd_sc_hd__nor2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6962_ clknet_leaf_88_core_clock _0223_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[15\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_214_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3321__S _0900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5102__A _1928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_76_core_clock_A clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_198_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5913_ _2681_ vssd1 vssd1 vccd1 vccd1 _2834_ sky130_fd_sc_hd__clkbuf_4
XFILLER_241_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6893_ clknet_leaf_76_core_clock _0154_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5844_ net201 vssd1 vssd1 vccd1 vccd1 _2791_ sky130_fd_sc_hd__buf_2
XANTENNA__4941__A _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4660__B _2081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5775_ _2681_ vssd1 vssd1 vccd1 vccd1 _2749_ sky130_fd_sc_hd__buf_2
XFILLER_158_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4152__S _1437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4726_ _2121_ immu_1.page_table\[6\]\[1\] _2123_ vssd1 vssd1 vccd1 vccd1 _2125_ sky130_fd_sc_hd__and3_1
XFILLER_147_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7445_ net74 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_1
X_4657_ _2072_ immu_1.page_table\[11\]\[10\] _2067_ vssd1 vssd1 vccd1 vccd1 _2080_
+ sky130_fd_sc_hd__and3_1
XFILLER_135_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3608_ _1190_ _1191_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__xor2_1
Xinput80 c0_sr_bus_addr[13] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
Xinput91 c0_sr_bus_addr[9] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_1
X_7376_ net301 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_2
XFILLER_162_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4588_ _1897_ vssd1 vssd1 vccd1 vccd1 _2038_ sky130_fd_sc_hd__buf_2
XFILLER_101_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6327_ _3069_ dmmu1.page_table\[3\]\[2\] _3077_ _3082_ vssd1 vssd1 vccd1 vccd1 _0498_
+ sky130_fd_sc_hd__a31o_1
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3539_ net153 dmmu1.long_off_reg\[3\] vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__or2_1
XFILLER_249_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3292__A _0869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6258_ _3026_ dmmu1.page_table\[5\]\[0\] _3038_ _3041_ vssd1 vssd1 vccd1 vccd1 _0470_
+ sky130_fd_sc_hd__a31o_1
XFILLER_249_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5655__A1 _2240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5209_ _2416_ dmmu0.page_table\[8\]\[7\] _2411_ vssd1 vssd1 vccd1 vccd1 _2420_ sky130_fd_sc_hd__and3_1
XFILLER_76_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6189_ _2998_ vssd1 vssd1 vccd1 vccd1 _2999_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4554__C _2004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6080__A1 _2932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3969__A1 _1479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3513__S0 _0896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4851__A _2084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3197__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input291_A ic0_mem_data[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input389_A inner_wb_i_dat[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4146__A1 _1411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5894__A1 _2239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6438__A3 _3135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7205__CLK clknet_leaf_28_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7402__A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6018__A _2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4082__B1 _1516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5857__A _2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3890_ net311 net365 _1390_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__mux2_1
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5560_ _2626_ vssd1 vssd1 vccd1 vccd1 _2627_ sky130_fd_sc_hd__clkbuf_4
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4511_ net207 vssd1 vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_11_core_clock clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_156_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5491_ _2590_ vssd1 vssd1 vccd1 vccd1 _2591_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5592__A _2640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7230_ clknet_leaf_23_core_clock _0491_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[4\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4442_ _1914_ _1930_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__nor2_4
XANTENNA__5885__A1 _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3824__B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7161_ clknet_leaf_9_core_clock _0422_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4373_ _1874_ _1875_ _1876_ _1806_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__a211o_1
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6112_ _2948_ dmmu1.page_table\[9\]\[7\] _2942_ _2953_ vssd1 vssd1 vccd1 vccd1 _0412_
+ sky130_fd_sc_hd__a31o_1
X_3324_ net17 vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__clkinv_4
X_7092_ clknet_leaf_35_core_clock _0353_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5637__A1 _2253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6043_ _2898_ dmmu1.page_table\[11\]\[6\] _2902_ _2911_ vssd1 vssd1 vccd1 vccd1 _0385_
+ sky130_fd_sc_hd__a31o_1
XFILLER_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3255_ net132 net27 _0847_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__mux2_2
XFILLER_273_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3840__A inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3186_ _0809_ _0810_ mem_dcache_arb.transfer_active vssd1 vssd1 vccd1 vccd1 net562
+ sky130_fd_sc_hd__a21oi_4
XFILLER_254_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4860__A2 _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4147__S _1453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ clknet_leaf_85_core_clock _0206_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[12\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_281_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3986__S _0811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5767__A _2736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_core_clock clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6876_ clknet_leaf_70_core_clock _0137_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5486__B _2577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5827_ _1946_ _2767_ _2779_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__a21o_1
XFILLER_210_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4376__A1 _1441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6872__CLK clknet_leaf_70_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5758_ _2235_ _2730_ _2739_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__a21o_1
XFILLER_6_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4709_ _2106_ immu_1.page_table\[9\]\[7\] _2103_ vssd1 vssd1 vccd1 vccd1 _2113_ sky130_fd_sc_hd__and3_1
XFILLER_5_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5689_ _2698_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7428_ net404 vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_1
XFILLER_118_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7228__CLK clknet_leaf_22_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4679__A2 _2083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7359_ net282 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_2
XANTENNA__3887__A0 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5340__A3 _2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5628__A1 _2245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4300__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4300__B2 _1411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input137_A c1_o_mem_data[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4057__S _0811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input304_A ic0_mem_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5800__A1 _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5396__B _2527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3925__A _1438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5867__A1 _2805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6020__B _2880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3878__A0 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5331__A3 _2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output523_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4756__A _2134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6745__CLK clknet_leaf_66_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput270 dcache_wb_o_dat[8] vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_8
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput281 ic0_mem_data[13] vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_1
XFILLER_236_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput292 ic0_mem_data[23] vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4842__A2 _2189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4991_ _2284_ immu_1.page_table\[15\]\[3\] _2282_ vssd1 vssd1 vccd1 vccd1 _2287_
+ sky130_fd_sc_hd__and3_1
XANTENNA__4055__B1 _1563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5587__A _2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4491__A _1968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6730_ clknet_leaf_66_core_clock _0800_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3942_ net368 vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__clkbuf_4
XFILLER_210_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6895__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6661_ clknet_leaf_80_core_clock _0731_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3873_ net250 _1393_ _1386_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__mux2_4
X_5612_ _2640_ dmmu0.page_table\[15\]\[1\] _2652_ vssd1 vssd1 vccd1 vccd1 _2654_ sky130_fd_sc_hd__and3_1
XANTENNA__5555__B1 _2625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6592_ clknet_leaf_44_core_clock _0662_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[9\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5543_ net85 net84 _2350_ vssd1 vssd1 vccd1 vccd1 _2621_ sky130_fd_sc_hd__or3_4
XFILLER_219_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5753__C _2732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5474_ net99 _2577_ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__and2_1
Xoutput700 net700 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[4] sky130_fd_sc_hd__buf_2
XFILLER_160_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5858__A1 _2618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7213_ clknet_leaf_23_core_clock _0474_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4425_ net82 net81 net80 net79 vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__or4_1
XFILLER_144_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3869__A0 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7144_ clknet_leaf_34_core_clock _0405_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_259_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4356_ immu_1.page_table\[8\]\[10\] immu_1.page_table\[9\]\[10\] _1439_ vssd1 vssd1
+ vccd1 vccd1 _1860_ sky130_fd_sc_hd__mux2_1
XFILLER_86_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3307_ _0896_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__buf_6
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7075_ clknet_leaf_10_core_clock _0336_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4287_ immu_0.page_table\[2\]\[9\] immu_0.page_table\[3\]\[9\] _1425_ vssd1 vssd1
+ vccd1 vccd1 _1792_ sky130_fd_sc_hd__mux2_1
XFILLER_274_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6026_ _2900_ vssd1 vssd1 vccd1 vccd1 _2901_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3238_ net118 net13 _0840_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__mux2_1
XFILLER_104_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6035__A1 _2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5497__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6928_ clknet_leaf_58_core_clock _0189_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5928__C _2832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6105__B _2944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6859_ clknet_leaf_72_core_clock _0120_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[7\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4349__A1 _1432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7050__CLK clknet_leaf_36_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3557__C1 _0957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3745__A _0839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6618__CLK clknet_leaf_53_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6121__A _1993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5849__A1 _2618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input254_A dcache_wb_adr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6768__CLK clknet_leaf_86_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4576__A _1999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4824__A2 _2172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4742__C _2123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5200__A _2400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6015__B _2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5854__B _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output640_A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5870__A _1989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4210_ immu_0.page_table\[2\]\[7\] immu_0.page_table\[3\]\[7\] net312 vssd1 vssd1
+ vccd1 vccd1 _1717_ sky130_fd_sc_hd__mux2_1
XANTENNA__3946__S0 _1437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5190_ _2217_ _2407_ vssd1 vssd1 vccd1 vccd1 _2408_ sky130_fd_sc_hd__nor2_1
XFILLER_79_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4141_ net7 immu_0.high_addr_off\[2\] vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__nor2_1
XFILLER_268_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4486__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6265__A1 _3042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4917__C _2221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4072_ immu_1.page_table\[8\]\[4\] immu_1.page_table\[9\]\[4\] immu_1.page_table\[10\]\[4\]
+ immu_1.page_table\[11\]\[4\] _1439_ _1581_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__mux4_2
XFILLER_256_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_15_core_clock_A clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_95_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4815__A2 _2172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4579__A1 _1996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4974_ _1981_ _2274_ _2277_ immu_1.page_table\[0\]\[6\] vssd1 vssd1 vccd1 vccd1 _0759_
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5748__C _2732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5110__A _1940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_1_core_clock clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__7073__CLK clknet_leaf_79_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3925_ _1438_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__buf_6
X_6713_ clknet_leaf_61_core_clock _0783_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[15\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_204_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6644_ clknet_leaf_56_core_clock _0714_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3856_ net231 _1381_ net664 vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__mux2_4
X_6575_ clknet_leaf_46_core_clock _0645_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3787_ _1344_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__clkbuf_1
XFILLER_164_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4160__S _1438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5526_ net98 _2609_ vssd1 vssd1 vccd1 vccd1 _2612_ sky130_fd_sc_hd__and2_1
XFILLER_117_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3284__B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6910__CLK clknet_leaf_76_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5457_ _2312_ _2559_ vssd1 vssd1 vccd1 vccd1 _2570_ sky130_fd_sc_hd__and2_1
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput530 net530 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[18] sky130_fd_sc_hd__buf_2
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5780__A _2749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput541 net541 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[6] sky130_fd_sc_hd__buf_2
Xoutput552 net552 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[15] sky130_fd_sc_hd__buf_2
XFILLER_160_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput563 net563 vssd1 vssd1 vccd1 vccd1 dcache_mem_sel[0] sky130_fd_sc_hd__buf_2
X_4408_ net664 _1579_ net388 vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__and3_1
XFILLER_278_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput574 net574 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[14] sky130_fd_sc_hd__buf_2
X_5388_ _2517_ immu_0.page_table\[7\]\[2\] _2525_ _2529_ vssd1 vssd1 vccd1 vccd1 _0112_
+ sky130_fd_sc_hd__a31o_1
Xoutput585 net585 vssd1 vssd1 vccd1 vccd1 ic0_clk sky130_fd_sc_hd__clkbuf_1
Xoutput596 net596 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[4] sky130_fd_sc_hd__buf_2
X_7127_ clknet_leaf_28_core_clock _0388_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[11\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4396__A _1895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4339_ _1478_ _1842_ _1535_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__o21ai_1
XFILLER_59_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4827__C _2174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7058_ clknet_leaf_80_core_clock _0319_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3609__A3 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6009_ _2803_ _2881_ vssd1 vssd1 vccd1 vccd1 _2890_ sky130_fd_sc_hd__and2_1
XFILLER_274_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6008__A1 _2884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7500__A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4019__B1 _1462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5658__C _2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5020__A _1935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4990__A1 _1972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input371_A ic1_wb_adr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6590__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input65_A c0_o_req_addr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3950__C1 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5690__A _2217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6495__A1 _1981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_6_0_core_clock_A clknet_2_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6247__A1 _3026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_6_core_clock_A clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_172_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7410__A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7096__CLK clknet_leaf_32_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4245__S _1480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5865__A _2561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3710_ _0905_ _1286_ _1288_ _1290_ net18 vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__o221a_1
X_4690_ _2100_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__clkbuf_4
XFILLER_201_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3641_ _1222_ _1223_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__nand2_1
XANTENNA__6933__CLK clknet_leaf_57_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5525__A3 _2607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4733__A1 _2012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6360_ _3101_ dmmu1.page_table\[2\]\[2\] _3096_ _3102_ vssd1 vssd1 vccd1 vccd1 _0511_
+ sky130_fd_sc_hd__a31o_1
X_3572_ dmmu1.page_table\[6\]\[9\] dmmu1.page_table\[7\]\[9\] _1146_ vssd1 vssd1 vccd1
+ vccd1 _1156_ sky130_fd_sc_hd__mux2_1
X_5311_ _1935_ _2482_ vssd1 vssd1 vccd1 vccd1 _2485_ sky130_fd_sc_hd__and2_1
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6291_ _3053_ dmmu1.page_table\[4\]\[0\] _3058_ _3061_ vssd1 vssd1 vccd1 vccd1 _0483_
+ sky130_fd_sc_hd__a31o_1
XFILLER_142_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5242_ _2444_ vssd1 vssd1 vccd1 vccd1 _2445_ sky130_fd_sc_hd__clkbuf_4
XFILLER_216_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3832__B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5173_ _2236_ _2390_ _2398_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__a21o_1
XANTENNA__3395__S1 _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4647__C _2068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4124_ _1440_ _1617_ _1618_ _1632_ _1360_ vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__o311a_2
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4249__B1 _1754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 c0_o_c_data_page vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_2
XFILLER_283_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4944__A _2262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4055_ _1553_ _1559_ _1563_ _1565_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__o22a_1
XFILLER_209_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4663__B _2081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4957_ _1985_ _2257_ _2269_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__a21o_1
XFILLER_196_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5775__A _2681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3908_ _1420_ _1421_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__nand2_1
XANTENNA__4972__A1 _1977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4888_ _2204_ dmmu0.page_table\[0\]\[0\] _2221_ vssd1 vssd1 vccd1 vccd1 _2222_ sky130_fd_sc_hd__and3_1
XFILLER_131_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5494__B _2589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3839_ _1372_ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_1
X_6627_ clknet_leaf_41_core_clock _0697_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3527__A2 _1088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6558_ clknet_leaf_50_core_clock _0628_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[12\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_83_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5509_ net103 _2593_ vssd1 vssd1 vccd1 vccd1 _2601_ sky130_fd_sc_hd__and2_1
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6489_ dmmu1.long_off_reg\[3\] _1974_ _3172_ vssd1 vssd1 vccd1 vccd1 _3176_ sky130_fd_sc_hd__mux2_1
XANTENNA__6477__A1 _1987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5015__A _1930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input217_A dcache_mem_o_data[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5204__A2 _2409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6956__CLK clknet_leaf_85_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3310__S1 _0902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6180__A3 _2981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7405__A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4748__B _2136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3377__S1 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output436_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4494__A3 _1964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4764__A _2134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4483__B _1961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3454__A1 dmmu0.page_table\[3\]\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5860_ _2801_ _2789_ vssd1 vssd1 vccd1 vccd1 _2802_ sky130_fd_sc_hd__and2_1
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4811_ _2006_ _2172_ _2176_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__a21o_1
XFILLER_33_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5791_ _2239_ _2748_ _2758_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__a21o_1
X_4742_ _2121_ immu_1.page_table\[6\]\[9\] _2123_ vssd1 vssd1 vccd1 vccd1 _2133_ sky130_fd_sc_hd__and3_1
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7461_ net400 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_1
X_4673_ _2010_ _2083_ _2091_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__a21o_1
XANTENNA__6203__B _3002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7111__CLK clknet_leaf_35_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6412_ net200 _3117_ vssd1 vssd1 vccd1 vccd1 _3132_ sky130_fd_sc_hd__and2_1
XANTENNA__4706__A1 _2014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3624_ _1205_ _1206_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__nand2_1
X_7392_ net362 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4004__A _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6343_ _2895_ _3078_ vssd1 vssd1 vccd1 vccd1 _3091_ sky130_fd_sc_hd__and2_1
X_3555_ _1138_ _1139_ _0917_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__mux2_2
XFILLER_115_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4939__A _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3843__A _1373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6459__A1 _1995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5761__C _2732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3390__B1 _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6274_ _2891_ _3040_ vssd1 vssd1 vccd1 vccd1 _3050_ sky130_fd_sc_hd__and2_1
XFILLER_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3486_ dmmu0.page_table\[12\]\[6\] dmmu0.page_table\[13\]\[6\] dmmu0.page_table\[14\]\[6\]
+ dmmu0.page_table\[15\]\[6\] _0900_ _0912_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__mux4_1
XFILLER_130_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5225_ _2081_ _2429_ vssd1 vssd1 vccd1 vccd1 _2430_ sky130_fd_sc_hd__nor2_2
XANTENNA__5131__A1 _2211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6829__CLK clknet_leaf_69_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5156_ _2253_ _2368_ _2387_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__a21o_1
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3989__S _1472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4107_ net111 immu_1.high_addr_off\[1\] vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__or2_1
XANTENNA__4674__A _2089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5087_ _2332_ immu_0.page_table\[12\]\[7\] _2336_ _2345_ vssd1 vssd1 vccd1 vccd1
+ _0804_ sky130_fd_sc_hd__a31o_1
XFILLER_217_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4038_ _1419_ _1548_ _1416_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__a21o_1
XANTENNA__6979__CLK clknet_leaf_57_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5001__C _2282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _2876_ vssd1 vssd1 vccd1 vccd1 _2877_ sky130_fd_sc_hd__clkbuf_2
XFILLER_12_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4945__A1 _1972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6113__B _2944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6162__A3 _2981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4849__A _1999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3753__A _1326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3381__B1 _0906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input167_A c1_o_req_addr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5122__A1 _2363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3191__C net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input334_A ic1_mem_data[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input28_A c0_o_mem_addr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4584__A _2017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3928__A net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7134__CLK clknet_leaf_13_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6023__B _2880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7284__CLK clknet_leaf_26_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3663__A _0901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3372__B1 _0855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3340_ dmmu1.page_table\[12\]\[1\] dmmu1.page_table\[13\]\[1\] _0857_ vssd1 vssd1
+ vccd1 vccd1 _0932_ sky130_fd_sc_hd__mux2_1
XANTENNA__5581__C _2634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A1 _2347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _0863_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__clkbuf_4
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _2297_ vssd1 vssd1 vccd1 vccd1 _2298_ sky130_fd_sc_hd__clkbuf_4
XFILLER_100_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6961_ clknet_leaf_88_core_clock _0222_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[15\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_226_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5102__B _2355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5912_ _2210_ _2830_ _2833_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__a21o_1
XFILLER_253_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_40_core_clock clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_179_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6892_ clknet_leaf_82_core_clock _0153_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[4\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_5843_ _2618_ dmmu1.page_table\[15\]\[0\] _2787_ _2790_ vssd1 vssd1 vccd1 vccd1 _0306_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__4941__B immu_1.page_table\[7\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3838__A _1363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4927__A1 _2249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6214__A _2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5774_ _2747_ vssd1 vssd1 vccd1 vccd1 _2748_ sky130_fd_sc_hd__clkbuf_4
XFILLER_166_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6392__A3 _3116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4725_ _1996_ _2120_ _2124_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__a21o_1
XFILLER_159_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4656_ _2023_ _2066_ _2079_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__a21o_1
X_7444_ net73 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_1
XFILLER_174_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3607_ _1130_ _1131_ _1129_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__a21bo_1
Xinput70 c0_o_req_addr[5] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__buf_2
XFILLER_135_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput81 c0_sr_bus_addr[14] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4669__A _1897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4587_ _2012_ _2030_ _2037_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__a21o_1
X_7375_ net300 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_2
Xinput92 c0_sr_bus_data_o[0] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_4
XANTENNA__6651__CLK clknet_leaf_38_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6326_ net202 _3079_ vssd1 vssd1 vccd1 vccd1 _3082_ sky130_fd_sc_hd__and2_1
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3538_ net153 dmmu1.long_off_reg\[3\] vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nand2_1
XFILLER_107_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6257_ _2879_ _3040_ vssd1 vssd1 vccd1 vccd1 _3041_ sky130_fd_sc_hd__and2_1
XFILLER_254_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3469_ _0957_ _1055_ _1056_ _0835_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__a31o_1
XFILLER_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5655__A2 _2669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5208_ _2240_ _2409_ _2419_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__a21o_1
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7007__CLK clknet_leaf_79_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6188_ _2919_ _2255_ vssd1 vssd1 vccd1 vccd1 _2998_ sky130_fd_sc_hd__or2_1
XFILLER_130_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5139_ _2233_ _2369_ _2378_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__a21o_1
XFILLER_111_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3512__S _0918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7157__CLK clknet_leaf_13_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3513__S1 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4851__B _2193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4343__S _1472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4918__A1 _2243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5666__C _2670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5591__A1 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5963__A _2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input284_A ic0_mem_data[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5894__A2 _2812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5203__A _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6018__B _2880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4082__A1 _1523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5857__B _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6034__A _2793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6374__A3 _3096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5582__A1 _2224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4510_ _1976_ dmmu1.page_table\[14\]\[6\] _1964_ _1982_ vssd1 vssd1 vccd1 vccd1 _0590_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__6674__CLK clknet_leaf_58_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3593__B1 _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5490_ _1929_ _2589_ vssd1 vssd1 vccd1 vccd1 _2590_ sky130_fd_sc_hd__or2_1
XFILLER_144_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5334__A1 _2489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4441_ _1929_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4489__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5885__A2 _2812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7160_ clknet_leaf_12_core_clock _0421_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4372_ _1807_ _1809_ vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__and2_1
XFILLER_208_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6111_ _2803_ _2944_ vssd1 vssd1 vccd1 vccd1 _2953_ sky130_fd_sc_hd__and2_1
X_3323_ _0909_ _0911_ _0915_ _0906_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__o211a_1
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7091_ clknet_leaf_2_core_clock _0352_ vssd1 vssd1 vccd1 vccd1 dmmu0.long_off_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6042_ _2801_ _2904_ vssd1 vssd1 vccd1 vccd1 _2911_ sky130_fd_sc_hd__and2_1
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3254_ _0850_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3648__A1 dmmu0.page_table\[3\]\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4845__B1 _2192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3185_ mem_dcache_arb.req1_pending net159 vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__nor2_4
XANTENNA__4655__C _2068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6944_ clknet_leaf_83_core_clock _0205_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4952__A _2262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6875_ clknet_leaf_71_core_clock _0136_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5826_ _2777_ dmmu0.page_table\[3\]\[8\] _2769_ vssd1 vssd1 vccd1 vccd1 _2779_ sky130_fd_sc_hd__and3_1
XFILLER_210_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4376__A2 _1864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5573__A1 _1948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5757_ _2736_ dmmu0.page_table\[4\]\[5\] _2732_ vssd1 vssd1 vccd1 vccd1 _2739_ sky130_fd_sc_hd__and3_1
XFILLER_210_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_opt_2_0_core_clock_A clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4708_ _2016_ _2101_ _2112_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_22_core_clock_A clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_175_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5688_ _2242_ immu_0.high_addr_off\[7\] _2690_ vssd1 vssd1 vccd1 vccd1 _2698_ sky130_fd_sc_hd__mux2_1
XFILLER_147_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4399__A _1897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7427_ net403 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5325__A1 _2489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4639_ _2006_ _2066_ _2070_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__a21o_1
XFILLER_118_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7358_ net281 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_2
XANTENNA__3887__A1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6309_ _2893_ _3060_ vssd1 vssd1 vccd1 vccd1 _3071_ sky130_fd_sc_hd__and2_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7289_ clknet_leaf_93_core_clock _0550_ vssd1 vssd1 vccd1 vccd1 mem_dcache_arb.req0_pending
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_277_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7503__A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5628__A2 _2650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_281_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4338__S _1480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6119__A _1991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3242__S _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3498__S0 _0891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5800__A2 _2747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4073__S _1439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6697__CLK clknet_leaf_42_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input95_A c0_sr_bus_data_o[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6108__A3 _2942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5316__A1 _2363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3422__S0 _0897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3878__A1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7413__A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput260 dcache_wb_o_dat[13] vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_1
XFILLER_283_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput271 dcache_wb_o_dat[9] vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_1
XFILLER_82_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput282 ic0_mem_data[14] vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_1
Xinput293 ic0_mem_data[24] vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5868__A _1987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4055__A1 _1553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4990_ _1972_ _2280_ _2286_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__a21o_1
XFILLER_251_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4491__B _1961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3941_ immu_1.page_table\[0\]\[0\] immu_1.page_table\[1\]\[0\] immu_1.page_table\[2\]\[0\]
+ immu_1.page_table\[3\]\[0\] _1453_ _1454_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__mux4_1
XFILLER_223_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6660_ clknet_leaf_7_core_clock _0730_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3872_ net320 net374 _1390_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__mux2_2
XFILLER_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5611_ _2211_ _2650_ _2653_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__a21o_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5555__A1 _2242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6591_ clknet_leaf_45_core_clock _0661_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[9\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5542_ _2618_ immu_0.page_table\[2\]\[10\] _2606_ _2620_ vssd1 vssd1 vccd1 vccd1
+ _0175_ sky130_fd_sc_hd__a31o_1
XFILLER_129_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5473_ _2576_ immu_0.page_table\[4\]\[3\] _2574_ _2580_ vssd1 vssd1 vccd1 vccd1 _0146_
+ sky130_fd_sc_hd__a31o_1
Xoutput701 net701 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[5] sky130_fd_sc_hd__buf_2
XANTENNA__5108__A _1937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4424_ _1912_ _1913_ vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__or2_4
X_7212_ clknet_leaf_16_core_clock _0473_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4012__A _1448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7143_ clknet_leaf_29_core_clock _0404_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[10\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_4355_ _1496_ _1858_ _1516_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_88_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_259_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3851__A _1373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3306_ net18 vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__buf_2
XFILLER_98_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7074_ clknet_leaf_79_core_clock _0335_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4286_ immu_0.page_table\[0\]\[9\] immu_0.page_table\[1\]\[9\] _1601_ vssd1 vssd1
+ vccd1 vccd1 _1791_ sky130_fd_sc_hd__mux2_1
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6025_ _2784_ _2064_ vssd1 vssd1 vccd1 vccd1 _2900_ sky130_fd_sc_hd__or2_1
X_3237_ _0841_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4158__S _1453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5778__A _2749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4682__A _2089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5497__B _2593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6927_ clknet_leaf_60_core_clock _0188_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_202_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3298__A _0857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6858_ clknet_leaf_69_core_clock _0119_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[7\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6338__A3 _3077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5809_ _2762_ dmmu0.page_table\[3\]\[0\] _2769_ vssd1 vssd1 vccd1 vccd1 _2770_ sky130_fd_sc_hd__and3_1
XFILLER_22_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6789_ clknet_leaf_3_core_clock _0050_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__dfxtp_2
XFILLER_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5018__A _1933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4857__A _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3761__A _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input247_A dcache_wb_adr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4576__B _2028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5077__A3 _2336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4285__A1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input10_A c0_o_instr_long_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5234__B1 _2434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_90_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5785__A1 _2229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6329__A3 _3077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5537__A1 _2603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3936__A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7408__A net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6712__CLK clknet_leaf_63_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output633_A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3946__S1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4140_ _1576_ _1610_ _1609_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__a21boi_2
XFILLER_95_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4071_ _1454_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__buf_4
XANTENNA__6862__CLK clknet_leaf_70_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4276__B2 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5598__A _2640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7218__CLK clknet_leaf_28_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4579__A2 _2030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4973_ _1979_ _2274_ _2277_ immu_1.page_table\[0\]\[5\] vssd1 vssd1 vccd1 vccd1 _0758_
+ sky130_fd_sc_hd__o22a_1
XFILLER_196_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5110__B _2355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6712_ clknet_leaf_63_core_clock _0782_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3924_ _1437_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__buf_6
XFILLER_149_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6643_ clknet_leaf_39_core_clock _0713_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3855_ net309 net363 _1360_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__mux2_2
XANTENNA__3846__A _1376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6222__A _3018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6574_ clknet_leaf_46_core_clock _0644_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3786_ net222 _0993_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__and2_1
XFILLER_192_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5525_ _2603_ immu_0.page_table\[2\]\[2\] _2607_ _2611_ vssd1 vssd1 vccd1 vccd1 _0167_
+ sky130_fd_sc_hd__a31o_1
XFILLER_117_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3284__C net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput520 net520 vssd1 vssd1 vccd1 vccd1 dcache_clk sky130_fd_sc_hd__clkbuf_1
X_5456_ _2562_ immu_0.page_table\[5\]\[8\] _2557_ _2569_ vssd1 vssd1 vccd1 vccd1 _0140_
+ sky130_fd_sc_hd__a31o_1
XFILLER_172_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput531 net531 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[19] sky130_fd_sc_hd__buf_2
XFILLER_59_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput542 net542 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[7] sky130_fd_sc_hd__buf_2
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput553 net553 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[1] sky130_fd_sc_hd__buf_2
X_4407_ _1903_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_1
Xoutput564 net564 vssd1 vssd1 vccd1 vccd1 dcache_mem_sel[1] sky130_fd_sc_hd__buf_2
Xoutput575 net575 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[15] sky130_fd_sc_hd__buf_2
X_5387_ _1933_ _2527_ vssd1 vssd1 vccd1 vccd1 _2529_ sky130_fd_sc_hd__and2_1
XFILLER_259_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput586 net586 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[0] sky130_fd_sc_hd__buf_2
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7126_ clknet_leaf_33_core_clock _0387_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[11\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput597 net597 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[5] sky130_fd_sc_hd__buf_2
X_4338_ immu_0.page_table\[10\]\[10\] immu_0.page_table\[11\]\[10\] _1480_ vssd1 vssd1
+ vccd1 vccd1 _1842_ sky130_fd_sc_hd__mux2_1
XFILLER_262_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input2_A c0_o_c_instr_long vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7057_ clknet_leaf_31_core_clock _0318_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[15\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_4269_ immu_1.page_table\[0\]\[8\] immu_1.page_table\[1\]\[8\] _1438_ vssd1 vssd1
+ vccd1 vccd1 _1775_ sky130_fd_sc_hd__mux2_1
XFILLER_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6008_ _2884_ dmmu1.page_table\[12\]\[6\] _2878_ _2889_ vssd1 vssd1 vccd1 vccd1 _0372_
+ sky130_fd_sc_hd__a31o_1
XFILLER_86_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4019__A1 _1457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5020__B _2302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4990__A2 _2280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input197_A c1_sr_bus_data_o[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5971__A _2561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input364_A ic1_wb_adr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5690__B _2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input58_A c0_o_req_active vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3466__C1 _1053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6307__A _2891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5211__A _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5758__A1 _2235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3233__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3640_ net50 dmmu0.long_off_reg\[5\] vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__or2_1
XANTENNA__6183__A1 _2994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6042__A _2801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3571_ _0869_ _1154_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__and2_1
XFILLER_174_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4733__A2 _2120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3941__A0 immu_1.page_table\[0\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5310_ _2363_ immu_0.page_table\[10\]\[2\] _2480_ _2484_ vssd1 vssd1 vccd1 vccd1
+ _0079_ sky130_fd_sc_hd__a31o_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6290_ _2879_ _3060_ vssd1 vssd1 vccd1 vccd1 _3061_ sky130_fd_sc_hd__and2_1
XFILLER_154_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5241_ _2443_ _2440_ vssd1 vssd1 vccd1 vccd1 _2444_ sky130_fd_sc_hd__or2_1
XFILLER_142_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4497__A1 _1939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5172_ _2384_ dmmu0.page_table\[9\]\[5\] _2392_ vssd1 vssd1 vccd1 vccd1 _2398_ sky130_fd_sc_hd__and3_1
XFILLER_275_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4123_ _1462_ _1625_ _1631_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__or3b_1
XFILLER_256_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4249__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4249__B2 _1411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 c0_o_c_instr_long vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_6
X_4054_ _1530_ _1564_ _1462_ _1457_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__a211o_1
XANTENNA__5997__A1 _2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7040__CLK clknet_leaf_12_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6608__CLK clknet_leaf_53_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5759__C _2732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3340__S _0857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5121__A _2314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5749__A1 _2223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4960__A _2262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4956_ _2262_ immu_1.page_table\[7\]\[8\] _2259_ vssd1 vssd1 vccd1 vccd1 _2269_ sky130_fd_sc_hd__and3_1
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3907_ immu_0.page_table\[14\]\[0\] immu_0.page_table\[15\]\[0\] _1408_ vssd1 vssd1
+ vccd1 vccd1 _1421_ sky130_fd_sc_hd__mux2_1
XANTENNA__4972__A2 _2274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4887_ _2220_ vssd1 vssd1 vccd1 vccd1 _2221_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__6174__A1 _2977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6626_ clknet_leaf_56_core_clock _0696_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3838_ _1363_ net270 vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__and2_1
XFILLER_118_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6557_ clknet_leaf_48_core_clock _0627_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[12\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3527__A3 _1095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5921__A1 _2232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3769_ _1334_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_1
XFILLER_257_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5508_ _2588_ immu_0.page_table\[3\]\[7\] _2591_ _2600_ vssd1 vssd1 vccd1 vccd1 _0161_
+ sky130_fd_sc_hd__a31o_1
XFILLER_145_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6488_ _3175_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_279_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6477__A2 _3157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5439_ net96 _2559_ vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__and2_1
XFILLER_126_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4488__A1 _1939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3515__S _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4200__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7109_ clknet_leaf_32_core_clock _0370_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5015__B _2296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5730__S _2720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5452__A3 _2557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4346__S _1407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6127__A _2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5031__A _2310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input112_A c1_o_instr_long_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4870__A _2204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3620__C1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4081__S _1439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5912__A1 _2210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5676__A0 _1928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7063__CLK clknet_leaf_10_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output429_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7421__A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5979__A1 _2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4256__S _1524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5579__C _2634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_core_clock clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6900__CLK clknet_leaf_75_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5876__A _2216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4810_ _2166_ immu_1.page_table\[2\]\[1\] _2174_ vssd1 vssd1 vccd1 vccd1 _2176_ sky130_fd_sc_hd__and3_1
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4780__A _2150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5790_ _2749_ dmmu0.page_table\[13\]\[6\] _2751_ vssd1 vssd1 vccd1 vccd1 _2758_ sky130_fd_sc_hd__and3_1
XFILLER_221_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4741_ _2021_ _2120_ _2132_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__a21o_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7460_ net399 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_1
X_4672_ _2089_ immu_1.page_table\[10\]\[3\] _2086_ vssd1 vssd1 vccd1 vccd1 _2091_
+ sky130_fd_sc_hd__and3_1
XFILLER_186_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6411_ _3128_ dmmu1.page_table\[1\]\[11\] _3115_ _3131_ vssd1 vssd1 vccd1 vccd1 _0533_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__4706__A2 _2101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3623_ net155 dmmu1.long_off_reg\[5\] vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__or2_1
X_7391_ net361 vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_1
XFILLER_227_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_27_core_clock_A clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_6342_ _3085_ dmmu1.page_table\[3\]\[9\] _3077_ _3090_ vssd1 vssd1 vccd1 vccd1 _0505_
+ sky130_fd_sc_hd__a31o_1
X_3554_ dmmu0.page_table\[8\]\[8\] dmmu0.page_table\[9\]\[8\] dmmu0.page_table\[10\]\[8\]
+ dmmu0.page_table\[11\]\[8\] _0896_ _0912_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__mux4_1
XFILLER_115_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6459__A2 _3157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6273_ _3042_ dmmu1.page_table\[5\]\[7\] _3038_ _3049_ vssd1 vssd1 vccd1 vccd1 _0477_
+ sky130_fd_sc_hd__a31o_1
X_3485_ _1070_ _1071_ _0918_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__mux2_1
XFILLER_115_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5116__A _2300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5224_ net196 net195 _1953_ _1956_ vssd1 vssd1 vccd1 vccd1 _2429_ sky130_fd_sc_hd__or4_2
XFILLER_130_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5131__A2 _2369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5155_ _2384_ dmmu0.page_table\[10\]\[12\] _2372_ vssd1 vssd1 vccd1 vccd1 _2387_
+ sky130_fd_sc_hd__and3_1
XFILLER_69_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4106_ net111 immu_1.high_addr_off\[1\] vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__nand2_1
XFILLER_272_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5086_ _1944_ _2338_ vssd1 vssd1 vccd1 vccd1 _2345_ sky130_fd_sc_hd__and2_1
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4037_ immu_0.page_table\[6\]\[3\] immu_0.page_table\[7\]\[3\] net312 vssd1 vssd1
+ vccd1 vccd1 _1548_ sky130_fd_sc_hd__mux2_1
XFILLER_244_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6580__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5786__A _2749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _2784_ _2045_ vssd1 vssd1 vccd1 vccd1 _2876_ sky130_fd_sc_hd__or2_1
XFILLER_241_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4939_ _2237_ immu_1.page_table\[7\]\[0\] _2259_ vssd1 vssd1 vccd1 vccd1 _2260_ sky130_fd_sc_hd__and3_1
XANTENNA__4945__A2 _2257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6147__A1 _1948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6609_ clknet_leaf_53_core_clock _0679_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7506__A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6410__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7086__CLK clknet_leaf_0_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4849__B _2193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5671__D _2212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4005__S0 _1453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5026__A _1942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4865__A _2105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input327_A ic0_wb_sel[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6923__CLK clknet_leaf_75_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5696__A _2682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6304__B _3060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6138__A1 _2235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7416__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6320__A _2784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3270_ _0860_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__clkbuf_4
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6310__A1 _3069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4775__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6960_ clknet_leaf_88_core_clock _0221_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[15\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4624__A1 _2021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5911_ _2819_ dmmu0.page_table\[5\]\[0\] _2832_ vssd1 vssd1 vccd1 vccd1 _2833_ sky130_fd_sc_hd__and3_1
XFILLER_241_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6891_ clknet_leaf_82_core_clock _0152_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[4\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5842_ _1995_ _2789_ vssd1 vssd1 vccd1 vccd1 _2790_ sky130_fd_sc_hd__and2_1
XFILLER_22_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4941__C _2259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4388__A0 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3838__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5773_ _2216_ _2351_ vssd1 vssd1 vccd1 vccd1 _2747_ sky130_fd_sc_hd__nor2_2
XFILLER_21_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4015__A _1442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4724_ _2121_ immu_1.page_table\[6\]\[0\] _2123_ vssd1 vssd1 vccd1 vccd1 _2124_ sky130_fd_sc_hd__and3_1
XFILLER_147_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7443_ net72 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_1
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4655_ _2072_ immu_1.page_table\[11\]\[9\] _2068_ vssd1 vssd1 vccd1 vccd1 _2079_
+ sky130_fd_sc_hd__and3_1
XFILLER_190_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3854__A _1380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3606_ _1188_ _1189_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__nand2_1
Xinput60 c0_o_req_addr[10] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_2
XFILLER_162_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput71 c0_o_req_addr[6] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_2
X_7374_ net298 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_2
X_4586_ _2017_ immu_1.page_table\[13\]\[4\] _2032_ vssd1 vssd1 vccd1 vccd1 _2037_
+ sky130_fd_sc_hd__and3_1
Xinput82 c0_sr_bus_addr[15] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_1
Xinput93 c0_sr_bus_data_o[10] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_2
XANTENNA__3363__A1 _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6325_ _3069_ dmmu1.page_table\[3\]\[1\] _3077_ _3081_ vssd1 vssd1 vccd1 vccd1 _0497_
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3537_ _0887_ _1115_ _1121_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__o21a_2
XFILLER_107_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6256_ _3039_ vssd1 vssd1 vccd1 vccd1 _3040_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__6301__A1 _3053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3468_ net45 dmmu0.long_off_reg\[0\] vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__or2_1
XANTENNA__6946__CLK clknet_leaf_81_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5207_ _2416_ dmmu0.page_table\[8\]\[6\] _2411_ vssd1 vssd1 vccd1 vccd1 _2419_ sky130_fd_sc_hd__and3_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6187_ _2994_ dmmu1.page_table\[8\]\[12\] _2980_ _2997_ vssd1 vssd1 vccd1 vccd1 _0443_
+ sky130_fd_sc_hd__a31o_1
XFILLER_191_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3399_ dmmu0.page_table\[8\]\[3\] dmmu0.page_table\[9\]\[3\] dmmu0.page_table\[10\]\[3\]
+ dmmu0.page_table\[11\]\[3\] _0898_ _0948_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__mux4_1
XFILLER_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5138_ _2371_ dmmu0.page_table\[10\]\[4\] _2373_ vssd1 vssd1 vccd1 vccd1 _2378_ sky130_fd_sc_hd__and3_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5069_ _1922_ _2334_ vssd1 vssd1 vccd1 vccd1 _2335_ sky130_fd_sc_hd__or2_1
XFILLER_270_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6080__A3 _2922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6405__A _1910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6368__A1 _3101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4918__A2 _2219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5591__A2 _2632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5963__B _2861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input277_A ic0_mem_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input40_A c0_o_mem_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4595__A _2038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4854__A1 _1995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3939__A _1437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6315__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7251__CLK clknet_leaf_19_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6034__B _2904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6819__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5582__A2 _2632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3593__A1 _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6480__B1_N _1899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3674__A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5592__C _2634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4440_ _1921_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__buf_4
XFILLER_7_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5334__A2 immu_0.page_table\[9\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6969__CLK clknet_leaf_86_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4371_ net116 immu_1.high_addr_off\[6\] vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__or2_1
XFILLER_208_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6110_ _2948_ dmmu1.page_table\[9\]\[6\] _2942_ _2952_ vssd1 vssd1 vccd1 vccd1 _0411_
+ sky130_fd_sc_hd__a31o_1
X_3322_ _0913_ _0914_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__or2_1
XFILLER_258_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7090_ clknet_leaf_2_core_clock _0351_ vssd1 vssd1 vccd1 vccd1 dmmu0.long_off_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6041_ _2898_ dmmu1.page_table\[11\]\[5\] _2902_ _2910_ vssd1 vssd1 vccd1 vccd1 _0384_
+ sky130_fd_sc_hd__a31o_1
XFILLER_85_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3253_ net131 net26 _0847_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__mux2_2
XANTENNA__4845__A1 _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3184_ mem_dcache_arb.req0_pending net54 vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__nor2_2
XFILLER_39_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6943_ clknet_leaf_85_core_clock _0204_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5270__A1 _2253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3849__A _1373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5767__C _2731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6874_ clknet_leaf_70_core_clock _0135_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6225__A _2879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5825_ _2242_ _2767_ _2778_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__a21o_1
XFILLER_210_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5756_ _2232_ _2730_ _2738_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__a21o_1
XFILLER_249_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4707_ _2106_ immu_1.page_table\[9\]\[6\] _2103_ vssd1 vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__and3_1
XFILLER_163_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5687_ _2697_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7426_ net402 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_1
X_4638_ _2054_ immu_1.page_table\[11\]\[1\] _2068_ vssd1 vssd1 vccd1 vccd1 _2070_
+ sky130_fd_sc_hd__and3_1
XFILLER_204_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7357_ net280 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_2
X_4569_ _1989_ vssd1 vssd1 vccd1 vccd1 _2025_ sky130_fd_sc_hd__buf_4
XFILLER_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6308_ _3069_ dmmu1.page_table\[4\]\[8\] _3058_ _3070_ vssd1 vssd1 vccd1 vccd1 _0491_
+ sky130_fd_sc_hd__a31o_1
XFILLER_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7288_ clknet_leaf_3_core_clock _0549_ vssd1 vssd1 vccd1 vccd1 mem_dcache_arb.req1_pending
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5089__A1 _2332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6239_ _3026_ dmmu1.page_table\[6\]\[6\] _3019_ _3029_ vssd1 vssd1 vccd1 vccd1 _0463_
+ sky130_fd_sc_hd__a31o_1
XFILLER_103_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7124__CLK clknet_leaf_34_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4297__C1 _1432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5304__A _1926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5261__A1 _2245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3498__S1 _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3759__A _1329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4354__S _1439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6135__A _2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3478__B _1064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5974__A _2801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input394_A inner_wb_i_dat[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input88_A c0_sr_bus_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5867__A3 _2787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3422__S1 _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4756__C _2140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput250 dcache_wb_adr[5] vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_4
XFILLER_236_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput261 dcache_wb_o_dat[14] vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_1
XFILLER_248_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput272 dcache_wb_sel[0] vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_4
Xinput283 ic0_mem_data[15] vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_1
Xinput294 ic0_mem_data[25] vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_1
XFILLER_263_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5868__B _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3940_ net367 vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__buf_4
XANTENNA__5587__C _2634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6641__CLK clknet_leaf_38_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3871_ _1392_ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__clkbuf_1
XFILLER_210_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5004__A1 _1987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5884__A _2777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5610_ _2640_ dmmu0.page_table\[15\]\[0\] _2652_ vssd1 vssd1 vccd1 vccd1 _2653_ sky130_fd_sc_hd__and3_1
X_6590_ clknet_leaf_45_core_clock _0660_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[9\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5555__A2 _2623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4212__C1 _1416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6791__CLK clknet_leaf_80_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5541_ net93 _2609_ vssd1 vssd1 vccd1 vccd1 _2620_ sky130_fd_sc_hd__and2_1
XFILLER_145_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5472_ net98 _2577_ vssd1 vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__and2_1
XFILLER_144_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput702 net702 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[6] sky130_fd_sc_hd__buf_2
X_7211_ clknet_leaf_16_core_clock _0472_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5108__B _2355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4423_ net84 net85 vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__or2b_1
XFILLER_132_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5858__A3 _2787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7147__CLK clknet_leaf_35_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7142_ clknet_leaf_29_core_clock _0403_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[10\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_4354_ immu_1.page_table\[12\]\[10\] immu_1.page_table\[13\]\[10\] _1439_ vssd1 vssd1
+ vccd1 vccd1 _1858_ sky130_fd_sc_hd__mux2_1
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3305_ _0897_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__buf_6
XFILLER_259_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7073_ clknet_leaf_79_core_clock _0334_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4285_ _1478_ _1787_ _1789_ _1479_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__o211a_1
XANTENNA__5124__A _2217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6024_ _2898_ dmmu1.page_table\[12\]\[12\] _2877_ _2899_ vssd1 vssd1 vccd1 vccd1
+ _0378_ sky130_fd_sc_hd__a31o_1
XANTENNA__7297__CLK clknet_leaf_43_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3236_ net162 net57 _0840_ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__mux2_1
XFILLER_239_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4963__A _1999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6035__A3 _2902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6926_ clknet_leaf_76_core_clock _0187_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6857_ clknet_leaf_69_core_clock _0118_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[7\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5794__A _2749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5808_ _2768_ vssd1 vssd1 vccd1 vccd1 _2769_ sky130_fd_sc_hd__buf_2
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6788_ clknet_leaf_2_core_clock _0049_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__dfxtp_2
XFILLER_210_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3557__A1 _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5739_ _2727_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7409_ net349 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5018__B _2302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5849__A3 _2787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6514__CLK clknet_leaf_36_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3253__S _0847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4809__A1 _1996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5034__A _2312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input142_A c1_o_mem_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4285__A2 _1787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5969__A _2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5234__A1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5234__B2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5785__A2 _2748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5200__C _2411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3428__S _0906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5209__A _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4113__A _1581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output459_A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7424__A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output626_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4070_ _1411_ _1575_ _1578_ _1579_ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__a211o_1
XANTENNA__6265__A3 _3038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5473__A1 _2576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3236__A0 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4972_ _1977_ _2274_ _2277_ immu_1.page_table\[0\]\[4\] vssd1 vssd1 vccd1 vccd1 _0757_
+ sky130_fd_sc_hd__o22a_1
XFILLER_251_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6711_ clknet_leaf_61_core_clock _0781_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3923_ net366 vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__buf_6
XFILLER_51_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6642_ clknet_leaf_56_core_clock _0712_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3854_ _1380_ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_1
X_6573_ clknet_leaf_46_core_clock _0643_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3785_ _1343_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__clkbuf_1
XFILLER_118_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5119__A _2312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4023__A _1534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5524_ net97 _2609_ vssd1 vssd1 vccd1 vccd1 _2611_ sky130_fd_sc_hd__and2_1
XANTENNA__6537__CLK clknet_leaf_44_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5455_ _2310_ _2559_ vssd1 vssd1 vccd1 vccd1 _2569_ sky130_fd_sc_hd__and2_1
XANTENNA__3284__D net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput510 net510 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[31] sky130_fd_sc_hd__buf_2
XANTENNA__4958__A _2262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput521 net521 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[0] sky130_fd_sc_hd__buf_2
XANTENNA__3862__A _0811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput532 net532 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[1] sky130_fd_sc_hd__buf_2
XANTENNA__5780__C _2751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput543 net543 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[8] sky130_fd_sc_hd__buf_2
X_4406_ net664 _1579_ net387 vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__and3_1
Xoutput554 net554 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[2] sky130_fd_sc_hd__buf_2
X_5386_ _2517_ immu_0.page_table\[7\]\[1\] _2525_ _2528_ vssd1 vssd1 vccd1 vccd1 _0111_
+ sky130_fd_sc_hd__a31o_1
Xoutput565 net565 vssd1 vssd1 vccd1 vccd1 dcache_mem_we sky130_fd_sc_hd__buf_2
Xoutput576 net576 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[1] sky130_fd_sc_hd__buf_2
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7125_ clknet_leaf_28_core_clock _0386_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput587 net587 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[10] sky130_fd_sc_hd__buf_2
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4337_ _1570_ _1840_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__nor2_1
Xoutput598 net598 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[6] sky130_fd_sc_hd__buf_2
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6687__CLK clknet_leaf_39_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7056_ clknet_leaf_31_core_clock _0317_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[15\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_259_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4268_ _1442_ _1773_ vssd1 vssd1 vccd1 vccd1 _1774_ sky130_fd_sc_hd__or2_1
X_6007_ _2801_ _2881_ vssd1 vssd1 vccd1 vccd1 _2889_ sky130_fd_sc_hd__and2_1
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4693__A _2089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3219_ _0830_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_1
XFILLER_27_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4199_ _1686_ _1687_ _1705_ _1462_ _1360_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__o221a_1
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6008__A3 _2878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5216__A1 _2249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_34_core_clock_A clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6909_ clknet_leaf_76_core_clock _0170_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4975__B1 _2277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5728__S _2720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3950__A1 _1439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4868__A _2204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input357_A ic1_mem_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4079__S _1524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6247__A3 _3018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3466__B1 _0929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_core_clock clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6307__B _3060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5758__A2 _2730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7419__A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6042__B _2904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3570_ dmmu1.page_table\[4\]\[9\] dmmu1.page_table\[5\]\[9\] _1146_ vssd1 vssd1 vccd1
+ vccd1 _1154_ sky130_fd_sc_hd__mux2_1
XFILLER_127_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4778__A _2084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _2215_ vssd1 vssd1 vccd1 vccd1 _2443_ sky130_fd_sc_hd__clkbuf_4
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5171_ _2233_ _2390_ _2397_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__a21o_1
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4122_ _1627_ _1629_ _1630_ _1456_ _1553_ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__a221o_1
XFILLER_256_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5446__A1 _2562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4053_ immu_1.page_table\[8\]\[3\] immu_1.page_table\[9\]\[3\] immu_1.page_table\[10\]\[3\]
+ immu_1.page_table\[11\]\[3\] _1438_ _1454_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__mux4_2
XFILLER_68_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput3 c0_o_c_instr_page vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_110_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5402__A _2312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4944__C _2259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5121__B _2355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4018__A _1451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5749__A2 _2730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4955_ _1983_ _2257_ _2268_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__a21o_1
XANTENNA__3857__A _1382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3906_ _1419_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__buf_4
XFILLER_177_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6233__A _2931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4886_ _2212_ _2215_ vssd1 vssd1 vccd1 vccd1 _2220_ sky130_fd_sc_hd__or2_1
XFILLER_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6625_ clknet_leaf_54_core_clock _0695_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[4\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3837_ _1371_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_1
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6556_ clknet_leaf_50_core_clock _0626_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5921__A2 _2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3768_ net139 net34 _0839_ vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__mux2_8
X_5507_ net102 _2593_ vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__and2_1
XFILLER_257_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6487_ dmmu1.long_off_reg\[2\] _1972_ _3172_ vssd1 vssd1 vccd1 vccd1 _3175_ sky130_fd_sc_hd__mux2_1
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3699_ _1280_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_1
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5438_ _1922_ _2555_ vssd1 vssd1 vccd1 vccd1 _2559_ sky130_fd_sc_hd__nor2_4
XFILLER_133_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5369_ _2517_ immu_0.page_table\[8\]\[5\] _2510_ _2518_ vssd1 vssd1 vccd1 vccd1 _0104_
+ sky130_fd_sc_hd__a31o_1
XFILLER_126_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7108_ clknet_leaf_37_core_clock _0369_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5437__A1 _2546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7039_ clknet_leaf_13_core_clock _0300_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6408__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3531__S _0857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6127__B dmmu0.page_table\[1\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5031__B _2302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input105_A c0_sr_bus_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6702__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3767__A _1333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6143__A _2681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5982__A _1989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6852__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5912__A2 _2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input70_A c0_o_req_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3706__S _1169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7208__CLK clknet_leaf_27_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5428__A1 _2546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3441__S _0857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4764__C _2140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5876__B _2539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6053__A _1991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4740_ _2121_ immu_1.page_table\[6\]\[8\] _2123_ vssd1 vssd1 vccd1 vccd1 _2132_ sky130_fd_sc_hd__and3_1
XFILLER_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4671_ _2008_ _2083_ _2090_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_3_2_0_core_clock_A clknet_2_1_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6410_ net199 _3117_ vssd1 vssd1 vccd1 vccd1 _3131_ sky130_fd_sc_hd__and2_1
XFILLER_174_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3622_ net155 dmmu1.long_off_reg\[5\] vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__nand2_1
X_7390_ net360 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_1
XFILLER_174_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6341_ _2893_ _3079_ vssd1 vssd1 vccd1 vccd1 _3090_ sky130_fd_sc_hd__and2_1
X_3553_ dmmu0.page_table\[12\]\[8\] dmmu0.page_table\[13\]\[8\] dmmu0.page_table\[14\]\[8\]
+ dmmu0.page_table\[15\]\[8\] _0896_ _0912_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__mux4_1
XANTENNA__3616__S net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4939__C _2259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6272_ _2803_ _3040_ vssd1 vssd1 vccd1 vccd1 _3049_ sky130_fd_sc_hd__and2_1
XANTENNA__4301__A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3484_ dmmu0.page_table\[0\]\[6\] dmmu0.page_table\[1\]\[6\] dmmu0.page_table\[2\]\[6\]
+ dmmu0.page_table\[3\]\[6\] _0900_ _0912_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__mux4_1
XFILLER_142_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5667__A1 _2251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5223_ _2367_ _2427_ vssd1 vssd1 vccd1 vccd1 _2428_ sky130_fd_sc_hd__and2b_1
XFILLER_102_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5154_ _2251_ _2368_ _2386_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__a21o_1
XFILLER_84_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4105_ _1411_ _1604_ _1608_ _1613_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__a31o_1
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5085_ _2332_ immu_0.page_table\[12\]\[6\] _2336_ _2344_ vssd1 vssd1 vccd1 vccd1
+ _0803_ sky130_fd_sc_hd__a31o_1
XFILLER_284_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4674__C _2086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5132__A _2371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4036_ immu_0.page_table\[4\]\[3\] immu_0.page_table\[5\]\[3\] _1472_ vssd1 vssd1
+ vccd1 vccd1 _1547_ sky130_fd_sc_hd__mux2_2
XANTENNA__6725__CLK clknet_leaf_62_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5987_ _2867_ dmmu1.page_table\[13\]\[12\] _2858_ _2875_ vssd1 vssd1 vccd1 vccd1
+ _0365_ sky130_fd_sc_hd__a31o_1
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3587__A _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6875__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4182__S _1443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4938_ _2258_ vssd1 vssd1 vccd1 vccd1 _2259_ sky130_fd_sc_hd__buf_2
XFILLER_268_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6147__A2 _2960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4869_ _1983_ _2195_ _2206_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__a21o_1
XFILLER_268_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6608_ clknet_leaf_53_core_clock _0678_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6539_ clknet_leaf_48_core_clock _0609_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6410__B _3117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5307__A _1928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4211__A _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4005__S1 _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5026__B _2302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4584__C _2032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5042__A _1922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input222_A dcache_mem_o_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6138__A2 _2960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7030__CLK clknet_leaf_7_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6320__B _2193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5217__A _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5649__A1 _2230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output441_A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7180__CLK clknet_leaf_29_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5113__A3 _2353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7432__A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4775__B net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4267__S _1453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6048__A _2561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6074__A1 _2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4624__A2 _2047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6898__CLK clknet_leaf_76_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5910_ _2831_ vssd1 vssd1 vccd1 vccd1 _2832_ sky130_fd_sc_hd__clkbuf_4
XFILLER_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6890_ clknet_leaf_82_core_clock _0151_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[4\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5841_ _2788_ vssd1 vssd1 vccd1 vccd1 _2789_ sky130_fd_sc_hd__clkbuf_4
XFILLER_234_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4572__B_N net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5772_ net95 _2729_ _2746_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__a21o_1
XFILLER_194_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4723_ _2122_ vssd1 vssd1 vccd1 vccd1 _2123_ sky130_fd_sc_hd__buf_2
XFILLER_238_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7442_ net71 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_1
X_4654_ _2021_ _2066_ _2078_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__a21o_1
XFILLER_238_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput50 c0_o_mem_high_addr[5] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
X_3605_ net49 dmmu0.long_off_reg\[4\] vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__or2_1
Xinput61 c0_o_req_addr[11] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_2
XFILLER_128_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7373_ net297 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_2
X_4585_ _2010_ _2030_ _2036_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__a21o_1
Xinput72 c0_o_req_addr[7] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_2
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5127__A _2370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput83 c0_sr_bus_addr[1] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_2
X_6324_ net201 _3079_ vssd1 vssd1 vccd1 vccd1 _3081_ sky130_fd_sc_hd__and2_1
Xinput94 c0_sr_bus_data_o[11] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_4
X_3536_ _1117_ _1119_ _1120_ _0881_ _0874_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__a221o_1
XANTENNA__3363__A2 _0947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6255_ _2784_ _2136_ vssd1 vssd1 vccd1 vccd1 _3039_ sky130_fd_sc_hd__nor2_1
XFILLER_130_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3467_ net45 dmmu0.long_off_reg\[0\] vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__nand2_1
XFILLER_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7342__A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5206_ _2236_ _2409_ _2418_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__a21o_1
X_6186_ _1993_ _2982_ vssd1 vssd1 vccd1 vccd1 _2997_ sky130_fd_sc_hd__and2_1
XFILLER_229_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3398_ _0921_ _0929_ _0987_ _0835_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__a31o_1
X_5137_ _2230_ _2369_ _2377_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__a21o_1
XFILLER_96_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5068_ net83 net76 _2295_ vssd1 vssd1 vccd1 vccd1 _2334_ sky130_fd_sc_hd__or3_4
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5812__A1 _2223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4019_ _1457_ _1529_ _1462_ _1530_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__a211o_1
XFILLER_272_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7053__CLK clknet_leaf_32_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5736__S _2720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6421__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5037__A _2314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input172_A c1_o_req_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4876__A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3780__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input33_A c0_o_mem_data[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4854__A2 _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6056__A1 _2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5203__C _2411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4067__B1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6315__B _3059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7427__A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5334__A3 _2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ net116 immu_1.high_addr_off\[6\] vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__nand2_1
XANTENNA__6570__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3321_ dmmu0.page_table\[12\]\[0\] dmmu0.page_table\[13\]\[0\] _0900_ vssd1 vssd1
+ vccd1 vccd1 _0914_ sky130_fd_sc_hd__mux2_1
XFILLER_171_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4786__A _2150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3690__A _0868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6295__A1 _3053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6040_ _2799_ _2904_ vssd1 vssd1 vccd1 vccd1 _2910_ sky130_fd_sc_hd__and2_1
X_3252_ _0849_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_1
XFILLER_100_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4845__A2 _2189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6047__A1 _2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6942_ clknet_leaf_85_core_clock _0203_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4952__C _2259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7076__CLK clknet_leaf_79_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3900__S0 _1407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6873_ clknet_leaf_70_core_clock _0134_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6225__B _3021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_core_clock_A clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_222_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4026__A _1535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5824_ _2777_ dmmu0.page_table\[3\]\[7\] _2769_ vssd1 vssd1 vccd1 vccd1 _2778_ sky130_fd_sc_hd__and3_1
XFILLER_249_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3569__C1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5755_ _2736_ dmmu0.page_table\[4\]\[4\] _2732_ vssd1 vssd1 vccd1 vccd1 _2738_ sky130_fd_sc_hd__and3_1
XFILLER_210_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4706_ _2014_ _2101_ _2111_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__a21o_1
XANTENNA__3584__A2 _1153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4781__A1 _1996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5686_ _2239_ immu_0.high_addr_off\[6\] _2690_ vssd1 vssd1 vccd1 vccd1 _2697_ sky130_fd_sc_hd__mux2_1
XFILLER_163_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6913__CLK clknet_leaf_79_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4637_ _1996_ _2066_ _2069_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__a21o_1
X_7425_ net401 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_1
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5325__A3 _2480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4568_ _2023_ _2002_ _2024_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__a21o_1
X_7356_ net279 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_2
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6307_ _2891_ _3060_ vssd1 vssd1 vccd1 vccd1 _3070_ sky130_fd_sc_hd__and2_1
X_3519_ net47 dmmu0.long_off_reg\[2\] vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__and2_1
XANTENNA__4696__A _2105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7287_ clknet_leaf_93_core_clock _0548_ vssd1 vssd1 vccd1 vccd1 mem_dcache_arb.select
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4499_ _1974_ _1970_ vssd1 vssd1 vccd1 vccd1 _1975_ sky130_fd_sc_hd__and2_1
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6238_ _2801_ _3021_ vssd1 vssd1 vccd1 vccd1 _3029_ sky130_fd_sc_hd__and2_1
XANTENNA__4297__B1 _1801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6169_ _2797_ _2983_ vssd1 vssd1 vccd1 vccd1 _2988_ sky130_fd_sc_hd__and2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6416__A _3134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5320__A _1944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5261__A2 _2442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5549__B1 _2625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5974__B _2861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4221__B1 _1410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3775__A _1337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4772__A1 _2023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input387_A inner_wb_ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6593__CLK clknet_leaf_59_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5316__A3 _2480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5990__A _2877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_41_core_clock_A clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_107_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6277__A1 _3042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput240 dcache_wb_adr[18] vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_2
XFILLER_236_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput251 dcache_wb_adr[6] vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_4
XANTENNA__7099__CLK clknet_leaf_32_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput262 dcache_wb_o_dat[15] vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_1
XFILLER_248_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput273 dcache_wb_sel[1] vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput284 ic0_mem_data[16] vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_1
Xinput295 ic0_mem_data[26] vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_1
XFILLER_263_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6326__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3870_ net249 _1391_ _1386_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__mux2_4
XANTENNA__5004__A2 _2280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5540_ _2618_ immu_0.page_table\[2\]\[9\] _2607_ _2619_ vssd1 vssd1 vccd1 vccd1 _0174_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__4763__A1 _2014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6061__A _1968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5471_ _2576_ immu_0.page_table\[4\]\[2\] _2574_ _2579_ vssd1 vssd1 vccd1 vccd1 _0145_
+ sky130_fd_sc_hd__a31o_1
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput703 net703 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[7] sky130_fd_sc_hd__buf_2
X_7210_ clknet_leaf_23_core_clock _0471_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4422_ net83 net76 vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__nand2_1
X_7141_ clknet_leaf_27_core_clock _0402_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[10\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4353_ _1523_ _1856_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__or2_1
XFILLER_235_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3304_ _0896_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__buf_6
X_7072_ clknet_leaf_79_core_clock _0333_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4284_ _1430_ _1788_ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__or2_1
X_6023_ _1993_ _2880_ vssd1 vssd1 vccd1 vccd1 _2899_ sky130_fd_sc_hd__and2_1
XANTENNA__5124__B _2367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3235_ _0839_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__buf_6
XFILLER_86_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4963__B _2272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5778__C _2751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6236__A _2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4682__C _2086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5140__A _2371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6440__A1 _1898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6925_ clknet_leaf_77_core_clock _0186_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_6856_ clknet_leaf_68_core_clock _0117_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5807_ _2443_ _2589_ vssd1 vssd1 vccd1 vccd1 _2768_ sky130_fd_sc_hd__or2_1
XFILLER_167_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3999_ immu_0.page_table\[12\]\[2\] immu_0.page_table\[13\]\[2\] _1472_ vssd1 vssd1
+ vccd1 vccd1 _1511_ sky130_fd_sc_hd__mux2_1
X_6787_ clknet_leaf_0_core_clock _0048_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[8\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4190__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3557__A2 _1137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5738_ immu_1.high_addr_off\[6\] _1981_ _2720_ vssd1 vssd1 vccd1 vccd1 _2727_ sky130_fd_sc_hd__mux2_1
XFILLER_129_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5669_ _2253_ _2668_ _2686_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__a21o_1
XFILLER_276_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7408_ net348 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__clkbuf_1
XFILLER_151_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4857__C _2197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5315__A _1940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5034__B _2302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4809__A2 _2172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6809__CLK clknet_leaf_86_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5969__B _2861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input135_A c1_o_mem_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_core_clock clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3493__B2 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_273_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4365__S _1439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6146__A _2971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5234__A2 _2433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input302_A ic0_mem_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5537__A3 _2607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5225__A _2081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7440__A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5598__C _2634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6422__A1 _3128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4971_ _1974_ _2274_ _2277_ immu_1.page_table\[0\]\[3\] vssd1 vssd1 vccd1 vccd1 _0756_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__5895__A _2819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6710_ clknet_leaf_63_core_clock _0780_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3922_ _1413_ _1418_ _1435_ _1411_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__o211ai_2
XFILLER_189_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3853_ _1373_ net262 vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__and2_4
X_6641_ clknet_leaf_38_core_clock _0711_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6572_ clknet_leaf_49_core_clock _0642_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3784_ net221 _0993_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__and2_1
XANTENNA__5119__B _2355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3944__C1 _1457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5523_ _2603_ immu_0.page_table\[2\]\[1\] _2607_ _2610_ vssd1 vssd1 vccd1 vccd1 _0166_
+ sky130_fd_sc_hd__a31o_1
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6489__A1 _1974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5454_ _2562_ immu_0.page_table\[5\]\[7\] _2557_ _2568_ vssd1 vssd1 vccd1 vccd1 _0139_
+ sky130_fd_sc_hd__a31o_1
XFILLER_133_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput500 net500 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[22] sky130_fd_sc_hd__buf_2
XFILLER_279_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7264__CLK clknet_leaf_19_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput511 net511 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[3] sky130_fd_sc_hd__buf_2
Xoutput522 net522 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[10] sky130_fd_sc_hd__buf_2
XFILLER_160_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4405_ _1902_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_1
Xoutput533 net533 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[20] sky130_fd_sc_hd__buf_2
Xoutput544 net544 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[9] sky130_fd_sc_hd__buf_2
X_5385_ net96 _2527_ vssd1 vssd1 vccd1 vccd1 _2528_ sky130_fd_sc_hd__and2_1
Xoutput555 net555 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[3] sky130_fd_sc_hd__buf_2
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput566 net566 vssd1 vssd1 vccd1 vccd1 dcache_rst sky130_fd_sc_hd__buf_2
Xoutput577 net577 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[2] sky130_fd_sc_hd__buf_2
X_7124_ clknet_leaf_34_core_clock _0385_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4336_ immu_0.page_table\[8\]\[10\] immu_0.page_table\[9\]\[10\] _1480_ vssd1 vssd1
+ vccd1 vccd1 _1840_ sky130_fd_sc_hd__mux2_1
XFILLER_5_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput588 net588 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[11] sky130_fd_sc_hd__buf_2
Xoutput599 net599 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[7] sky130_fd_sc_hd__buf_2
XFILLER_99_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7055_ clknet_leaf_30_core_clock _0316_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[15\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_247_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4267_ immu_1.page_table\[4\]\[8\] immu_1.page_table\[5\]\[8\] _1453_ vssd1 vssd1
+ vccd1 vccd1 _1773_ sky130_fd_sc_hd__mux2_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6006_ _2884_ dmmu1.page_table\[12\]\[5\] _2878_ _2888_ vssd1 vssd1 vccd1 vccd1 _0371_
+ sky130_fd_sc_hd__a31o_1
X_3218_ net229 _0824_ vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__and2_1
X_4198_ _1553_ _1691_ _1695_ _1704_ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__o31ai_1
XFILLER_255_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4185__S _1493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6413__A1 _3128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6908_ clknet_leaf_75_core_clock _0169_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4975__A1 _1983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6839_ clknet_leaf_68_core_clock _0100_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4188__C1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4727__A1 _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3950__A2 _1441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5152__A1 _2249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4360__C1 _1457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input252_A dcache_wb_adr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4884__A _2212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6781__CLK clknet_leaf_86_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6404__A1 _3112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5211__C _2411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7137__CLK clknet_leaf_34_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6183__A3 _2980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7287__CLK clknet_leaf_93_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7435__A clknet_opt_1_0_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4778__B _2153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5143__A1 _2240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4497__A3 _1964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5170_ _2384_ dmmu0.page_table\[9\]\[4\] _2392_ vssd1 vssd1 vccd1 vccd1 _2397_ sky130_fd_sc_hd__and3_1
XANTENNA__4351__C1 _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4121_ immu_1.page_table\[4\]\[5\] immu_1.page_table\[5\]\[5\] immu_1.page_table\[6\]\[5\]
+ immu_1.page_table\[7\]\[5\] _1493_ _1442_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__mux4_1
XFILLER_268_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6485__S _3172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4794__A _2150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4052_ _1523_ _1560_ _1562_ _1456_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__o211a_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 c0_o_icache_flush vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_2
XFILLER_49_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5997__A3 _2878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5402__B _2527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3203__A net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4957__A1 _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4954_ _2262_ immu_1.page_table\[7\]\[7\] _2259_ vssd1 vssd1 vccd1 vccd1 _2268_ sky130_fd_sc_hd__and3_1
XFILLER_196_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6504__CLK clknet_leaf_59_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3905_ net313 vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__buf_4
XFILLER_177_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4885_ _2218_ vssd1 vssd1 vccd1 vccd1 _2219_ sky130_fd_sc_hd__buf_4
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6624_ clknet_leaf_54_core_clock _0694_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[4\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3836_ _1363_ net269 vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__and2_1
XFILLER_137_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6174__A3 _2981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6555_ clknet_leaf_50_core_clock _0625_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3767_ _1333_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_1
XFILLER_192_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5506_ _2588_ immu_0.page_table\[3\]\[6\] _2591_ _2599_ vssd1 vssd1 vccd1 vccd1 _0160_
+ sky130_fd_sc_hd__a31o_1
XFILLER_3_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3698_ _1254_ _1279_ _0835_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__mux2_4
X_6486_ _3174_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5437_ _2546_ immu_0.page_table\[5\]\[0\] _2557_ _2558_ vssd1 vssd1 vccd1 vccd1 _0132_
+ sky130_fd_sc_hd__a31o_1
XFILLER_279_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4488__A3 _1964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5368_ _1940_ _2512_ vssd1 vssd1 vccd1 vccd1 _2518_ sky130_fd_sc_hd__and2_1
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7107_ clknet_leaf_36_core_clock _0368_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4319_ _1584_ _1823_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__or2_1
XFILLER_141_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5299_ _2251_ _2461_ _2477_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__a21o_1
X_7038_ clknet_leaf_9_core_clock _0299_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6408__B _3117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6127__C _2962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4870__C _2197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3259__S _0847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5373__A1 _2517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input63_A c0_o_req_addr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5503__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5979__A3 _2859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6527__CLK clknet_leaf_42_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4780__C _2157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3611__A1 _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6677__CLK clknet_leaf_56_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4670_ _2089_ immu_1.page_table\[10\]\[2\] _2086_ vssd1 vssd1 vccd1 vccd1 _2090_
+ sky130_fd_sc_hd__and3_1
XFILLER_119_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3621_ net123 _1197_ _1203_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__o21a_2
XANTENNA__5364__A1 _2503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3693__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6340_ _3085_ dmmu1.page_table\[3\]\[8\] _3077_ _3089_ vssd1 vssd1 vccd1 vccd1 _0504_
+ sky130_fd_sc_hd__a31o_1
X_3552_ _1135_ _1136_ _0918_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__mux2_1
XFILLER_174_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6271_ _3042_ dmmu1.page_table\[5\]\[6\] _3038_ _3048_ vssd1 vssd1 vccd1 vccd1 _0476_
+ sky130_fd_sc_hd__a31o_1
X_3483_ dmmu0.page_table\[4\]\[6\] dmmu0.page_table\[5\]\[6\] dmmu0.page_table\[6\]\[6\]
+ dmmu0.page_table\[7\]\[6\] _0900_ _0902_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__mux4_1
X_5222_ _1919_ _2426_ vssd1 vssd1 vccd1 vccd1 _2427_ sky130_fd_sc_hd__nor2_1
XANTENNA__4324__C1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5153_ _2384_ dmmu0.page_table\[10\]\[11\] _2372_ vssd1 vssd1 vccd1 vccd1 _2386_
+ sky130_fd_sc_hd__and3_1
XFILLER_229_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7302__CLK clknet_leaf_62_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4104_ net2 _1611_ _1612_ _1360_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__a31o_2
XFILLER_229_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5084_ _1942_ _2338_ vssd1 vssd1 vccd1 vccd1 _2344_ sky130_fd_sc_hd__and2_1
XFILLER_284_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4035_ _1419_ _1543_ _1545_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__a21o_1
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4029__A _1419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3868__A _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6244__A _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5786__C _2751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ _1993_ _2860_ vssd1 vssd1 vccd1 vccd1 _2875_ sky130_fd_sc_hd__and2_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4937_ _2084_ _2255_ vssd1 vssd1 vccd1 vccd1 _2258_ sky130_fd_sc_hd__or2_1
XANTENNA__3602__A1 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4868_ _2204_ immu_1.page_table\[3\]\[7\] _2197_ vssd1 vssd1 vccd1 vccd1 _2206_ sky130_fd_sc_hd__and3_1
XFILLER_227_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6607_ clknet_leaf_53_core_clock _0677_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4699__A _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3819_ net274 _1361_ net664 vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__mux2_4
X_4799_ _2166_ immu_1.page_table\[4\]\[9\] _2157_ vssd1 vssd1 vccd1 vccd1 _2168_ sky130_fd_sc_hd__and3_1
X_6538_ clknet_leaf_48_core_clock _0608_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5107__A1 _2347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5307__B _2482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6469_ _1979_ _3157_ _3165_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__a21o_1
XFILLER_137_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_46_core_clock_A clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_161_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6419__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5042__B _2318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4094__A1 _1535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input215_A dcache_mem_o_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6154__A _2931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5696__C _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5993__A _2880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4402__A _1898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5649__A2 _2669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__A3 _3058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output434_A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3452__S _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3688__A _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4717__B_N net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4283__S _1425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5840_ _1968_ _2278_ vssd1 vssd1 vccd1 vccd1 _2788_ sky130_fd_sc_hd__nor2_1
XFILLER_207_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5771_ _2736_ dmmu0.page_table\[4\]\[12\] _2731_ vssd1 vssd1 vccd1 vccd1 _2746_ sky130_fd_sc_hd__and3_1
XFILLER_222_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4722_ _2084_ _2118_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__or2_1
XFILLER_159_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7441_ net70 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_1
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4653_ _2072_ immu_1.page_table\[11\]\[8\] _2068_ vssd1 vssd1 vccd1 vccd1 _2078_
+ sky130_fd_sc_hd__and3_1
XFILLER_147_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput40 c0_o_mem_data[5] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4312__A _1581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3604_ net49 dmmu0.long_off_reg\[4\] vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__nand2_1
XFILLER_238_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput51 c0_o_mem_high_addr[6] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
X_7372_ net296 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_2
X_4584_ _2017_ immu_1.page_table\[13\]\[3\] _2032_ vssd1 vssd1 vccd1 vccd1 _2036_
+ sky130_fd_sc_hd__and3_1
Xinput62 c0_o_req_addr[12] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_2
Xinput73 c0_o_req_addr[8] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_2
XFILLER_128_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput84 c0_sr_bus_addr[2] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_2
X_6323_ _3069_ dmmu1.page_table\[3\]\[0\] _3077_ _3080_ vssd1 vssd1 vccd1 vccd1 _0496_
+ sky130_fd_sc_hd__a31o_1
Xinput95 c0_sr_bus_data_o[12] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_4
X_3535_ dmmu1.page_table\[8\]\[8\] dmmu1.page_table\[9\]\[8\] dmmu1.page_table\[10\]\[8\]
+ dmmu1.page_table\[11\]\[8\] _0865_ _0863_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__mux4_1
XANTENNA__4031__B _1410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6254_ _3037_ vssd1 vssd1 vccd1 vccd1 _3038_ sky130_fd_sc_hd__buf_4
X_3466_ _1039_ _1044_ _0929_ _1053_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__o211a_1
XFILLER_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6301__A3 _3058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5205_ _2416_ dmmu0.page_table\[8\]\[5\] _2411_ vssd1 vssd1 vccd1 vccd1 _2418_ sky130_fd_sc_hd__and3_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6185_ _2994_ dmmu1.page_table\[8\]\[11\] _2980_ _2996_ vssd1 vssd1 vccd1 vccd1 _0442_
+ sky130_fd_sc_hd__a31o_1
X_3397_ _0985_ _0986_ _0906_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__mux2_1
XFILLER_130_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5136_ _2371_ dmmu0.page_table\[10\]\[3\] _2373_ vssd1 vssd1 vccd1 vccd1 _2377_ sky130_fd_sc_hd__and3_1
XFILLER_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4982__A _2084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5067_ _2332_ immu_0.page_table\[14\]\[10\] _2319_ _2333_ vssd1 vssd1 vccd1 vccd1
+ _0796_ sky130_fd_sc_hd__a31o_1
XFILLER_229_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6842__CLK clknet_leaf_69_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4018_ _1451_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__buf_4
XFILLER_177_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3598__A _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4193__S _1443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6368__A3 _3096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6992__CLK clknet_leaf_9_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5969_ _2797_ _2861_ vssd1 vssd1 vccd1 vccd1 _2866_ sky130_fd_sc_hd__and2_1
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6421__B _3137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5037__B _2302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input165_A c1_o_req_addr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4839__B1 _2192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3780__B _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5500__A1 _2588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput400 inner_wb_i_dat[5] vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_8
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4595__C _2032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5053__A _1937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input332_A ic1_mem_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5988__A _2784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input26_A c0_o_mem_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4892__A _2204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4067__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5567__A1 _2229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3578__B1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7443__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3750__A0 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3320_ _0912_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__buf_4
XFILLER_98_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3251_ net130 net25 _0847_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__mux2_2
XFILLER_86_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6865__CLK clknet_leaf_70_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3502__B1 _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6493__S _3172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6452__C1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6941_ clknet_leaf_82_core_clock _0202_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_240_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3900__S1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6872_ clknet_leaf_70_core_clock _0133_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_234_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5558__A1 _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5823_ _2681_ vssd1 vssd1 vccd1 vccd1 _2777_ sky130_fd_sc_hd__clkbuf_4
XFILLER_179_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5754_ _2229_ _2730_ _2737_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__a21o_1
XFILLER_249_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4705_ _2106_ immu_1.page_table\[9\]\[5\] _2103_ vssd1 vssd1 vccd1 vccd1 _2111_ sky130_fd_sc_hd__and3_1
XANTENNA__3584__A3 _1162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4781__A2 _2155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5685_ _2696_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5138__A _2371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4042__A net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7424_ net400 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_1
X_4636_ _2054_ immu_1.page_table\[11\]\[0\] _2068_ vssd1 vssd1 vccd1 vccd1 _2069_
+ sky130_fd_sc_hd__and3_1
XFILLER_135_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7355_ net278 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_2
XANTENNA__5730__A1 _1972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4567_ _2017_ immu_1.page_table\[14\]\[9\] _2004_ vssd1 vssd1 vccd1 vccd1 _2024_
+ sky130_fd_sc_hd__and3_1
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3741__A0 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6306_ _2931_ vssd1 vssd1 vccd1 vccd1 _3069_ sky130_fd_sc_hd__buf_4
X_3518_ _0818_ _0928_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__nor2_1
X_7286_ clknet_leaf_26_core_clock _0547_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_4498_ net203 vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__buf_6
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5089__A3 _2336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6237_ _3026_ dmmu1.page_table\[6\]\[5\] _3019_ _3028_ vssd1 vssd1 vccd1 vccd1 _0462_
+ sky130_fd_sc_hd__a31o_1
XFILLER_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3449_ dmmu0.page_table\[4\]\[5\] dmmu0.page_table\[5\]\[5\] _0910_ vssd1 vssd1 vccd1
+ vccd1 _1037_ sky130_fd_sc_hd__mux2_1
XANTENNA__4297__A1 _1424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6168_ _2977_ dmmu1.page_table\[8\]\[3\] _2981_ _2987_ vssd1 vssd1 vccd1 vccd1 _0434_
+ sky130_fd_sc_hd__a31o_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _2312_ _2355_ vssd1 vssd1 vccd1 vccd1 _2365_ sky130_fd_sc_hd__and2_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6099_ _2932_ dmmu1.page_table\[9\]\[1\] _2942_ _2946_ vssd1 vssd1 vccd1 vccd1 _0406_
+ sky130_fd_sc_hd__a31o_1
XFILLER_27_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5797__A1 _1948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5320__B _2482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6135__C _2962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5549__A1 _2223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7170__CLK clknet_leaf_35_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6738__CLK clknet_leaf_66_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4772__A2 _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input282_A ic0_mem_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5721__A1 _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput230 dcache_wb_4_burst vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_1
XFILLER_283_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput241 dcache_wb_adr[19] vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
Xinput252 dcache_wb_adr[7] vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_4
XFILLER_276_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput263 dcache_wb_o_dat[1] vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_6
Xinput274 dcache_wb_stb vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_2
XANTENNA__3730__S _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5511__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput285 ic0_mem_data[17] vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput296 ic0_mem_data[27] vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_1
XFILLER_84_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_89_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__6326__B _3079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4460__A1 _1939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3966__A _1432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7438__A net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5884__C _2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4212__A1 _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6061__B _2081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4763__A2 _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5470_ net97 _2577_ vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__and2_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4421_ _1910_ vssd1 vssd1 vccd1 vccd1 _1911_ sky130_fd_sc_hd__buf_8
Xoutput704 net704 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[8] sky130_fd_sc_hd__buf_2
XANTENNA__4797__A _2166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5712__A1 _2245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7140_ clknet_leaf_29_core_clock _0401_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[10\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_4352_ immu_1.page_table\[14\]\[10\] immu_1.page_table\[15\]\[10\] _1524_ vssd1 vssd1
+ vccd1 vccd1 _1856_ sky130_fd_sc_hd__mux2_1
XFILLER_259_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3303_ _0895_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__buf_6
X_4283_ immu_0.page_table\[4\]\[9\] immu_0.page_table\[5\]\[9\] _1425_ vssd1 vssd1
+ vccd1 vccd1 _1788_ sky130_fd_sc_hd__mux2_1
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7071_ clknet_leaf_79_core_clock _0332_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3206__A _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3234_ _0838_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__clkbuf_8
X_6022_ _2561_ vssd1 vssd1 vccd1 vccd1 _2898_ sky130_fd_sc_hd__buf_4
XFILLER_246_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5421__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5779__A1 _2210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6236__B _3021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7193__CLK clknet_leaf_29_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6924_ clknet_leaf_58_core_clock _0185_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6855_ clknet_leaf_69_core_clock _0116_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5794__C _2751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5806_ _2766_ vssd1 vssd1 vccd1 vccd1 _2767_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__6252__A _2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6786_ clknet_leaf_0_core_clock _0047_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[8\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3998_ immu_0.page_table\[14\]\[2\] immu_0.page_table\[15\]\[2\] _1408_ vssd1 vssd1
+ vccd1 vccd1 _1510_ sky130_fd_sc_hd__mux2_1
XFILLER_200_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5737_ _2726_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5668_ _2682_ dmmu0.page_table\[11\]\[12\] _2670_ vssd1 vssd1 vccd1 vccd1 _2686_
+ sky130_fd_sc_hd__and3_1
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7407_ net347 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_1
X_4619_ _2054_ immu_1.page_table\[12\]\[6\] _2049_ vssd1 vssd1 vccd1 vccd1 _2057_
+ sky130_fd_sc_hd__and3_1
XANTENNA__5703__A1 _2233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4062__S0 _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5599_ _2247_ _2632_ _2645_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__a21o_1
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5315__B _2482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7269_ clknet_leaf_24_core_clock _0530_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6427__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input128_A c1_o_mem_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6560__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3786__A net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input93_A c0_sr_bus_data_o[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5942__A1 _1928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5209__C _2411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4053__S0 _1438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4410__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7066__CLK clknet_leaf_10_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5940__S _2848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5473__A3 _2574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4681__A1 _2019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5241__A _2443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6903__CLK clknet_leaf_76_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _1972_ _2274_ _2277_ immu_1.page_table\[0\]\[2\] vssd1 vssd1 vccd1 vccd1 _0755_
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3921_ _1422_ _1427_ _1429_ _1433_ _1434_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__a221o_1
XFILLER_189_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6640_ clknet_leaf_57_core_clock _0710_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3852_ _1379_ vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_1
XFILLER_204_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6571_ clknet_leaf_46_core_clock _0641_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5933__A1 _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3783_ _1342_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_1
XFILLER_192_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5522_ net96 _2609_ vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__and2_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5453_ net102 _2559_ vssd1 vssd1 vccd1 vccd1 _2568_ sky130_fd_sc_hd__and2_1
XFILLER_246_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput501 net501 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[23] sky130_fd_sc_hd__buf_2
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4958__C _2259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5416__A _2300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput512 net512 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[4] sky130_fd_sc_hd__buf_2
Xoutput523 net523 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[11] sky130_fd_sc_hd__buf_2
X_4404_ icore_sregs.c1_disable net384 vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__or2_1
Xoutput534 net534 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[21] sky130_fd_sc_hd__buf_2
Xoutput545 net545 vssd1 vssd1 vccd1 vccd1 dcache_mem_cache_enable sky130_fd_sc_hd__buf_2
X_5384_ _1930_ _2440_ vssd1 vssd1 vccd1 vccd1 _2527_ sky130_fd_sc_hd__nor2_4
Xoutput556 net556 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[4] sky130_fd_sc_hd__buf_2
Xoutput567 net567 vssd1 vssd1 vccd1 vccd1 dcache_wb_ack sky130_fd_sc_hd__buf_2
XFILLER_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7123_ clknet_leaf_13_core_clock _0384_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_259_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput578 net578 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[3] sky130_fd_sc_hd__buf_2
X_4335_ _1420_ _1838_ _1432_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__o21ai_1
XFILLER_259_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput589 net589 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[12] sky130_fd_sc_hd__buf_2
XFILLER_259_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7054_ clknet_leaf_31_core_clock _0315_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[15\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6110__A1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4266_ _1584_ _1771_ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__or2_1
XFILLER_247_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6005_ _2799_ _2881_ vssd1 vssd1 vccd1 vccd1 _2888_ sky130_fd_sc_hd__and2_1
X_3217_ _0829_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4693__C _2103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4197_ _1457_ _1699_ _1703_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__or3_2
XFILLER_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5151__A _2384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6583__CLK clknet_leaf_42_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_255_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ clknet_leaf_82_core_clock _0168_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_270_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3632__C1 _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4975__A2 _2274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6838_ clknet_leaf_68_core_clock _0099_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4727__A2 _2120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6769_ clknet_leaf_90_core_clock _0030_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7089__CLK clknet_leaf_2_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5688__A0 _2242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4868__C _2197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5326__A _2314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6101__A1 _2932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input245_A dcache_wb_adr[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4884__B _2217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6926__CLK clknet_leaf_76_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5061__A _2310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5996__A _2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_53_core_clock_A clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6168__A1 _2977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5915__A1 _2223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6340__A1 _3085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5143__A2 _2369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4351__B1 _1854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output631_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7451__A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4120_ _1584_ _1628_ _1451_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__o21a_1
XFILLER_1_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5446__A3 _2557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4286__S _1601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4051_ _1442_ _1561_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__or2_1
XANTENNA__6067__A _2793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4654__A1 _2021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 c0_o_instr_long_addr[0] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_4
XFILLER_237_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3203__B _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4957__A2 _2257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4953_ _1981_ _2257_ _2267_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__a21o_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3904_ _1417_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__inv_2
X_4884_ _2212_ _2217_ vssd1 vssd1 vccd1 vccd1 _2218_ sky130_fd_sc_hd__nor2_1
XFILLER_220_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6623_ clknet_leaf_54_core_clock _0693_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[4\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3835_ _1370_ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5906__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6554_ clknet_leaf_50_core_clock _0624_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_257_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3766_ net138 net33 _0839_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__mux2_4
X_5505_ net101 _2593_ vssd1 vssd1 vccd1 vccd1 _2599_ sky130_fd_sc_hd__and2_1
XFILLER_173_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6485_ dmmu1.long_off_reg\[1\] _1967_ _3172_ vssd1 vssd1 vccd1 vccd1 _3174_ sky130_fd_sc_hd__mux2_1
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4017__S0 _1438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3697_ _0879_ _1258_ _1259_ _1278_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__o31ai_4
XANTENNA__5146__A _2371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5436_ _1925_ _2556_ vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__nor2_1
XFILLER_133_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6331__A1 _3069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6949__CLK clknet_leaf_7_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5367_ _2300_ vssd1 vssd1 vccd1 vccd1 _2517_ sky130_fd_sc_hd__clkbuf_4
XFILLER_273_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4893__A1 _2224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7106_ clknet_leaf_32_core_clock _0367_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4318_ immu_1.page_table\[2\]\[9\] immu_1.page_table\[3\]\[9\] _1493_ vssd1 vssd1
+ vccd1 vccd1 _1823_ sky130_fd_sc_hd__mux2_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5298_ _2473_ dmmu0.page_table\[14\]\[11\] _2463_ vssd1 vssd1 vccd1 vccd1 _2477_
+ sky130_fd_sc_hd__and3_1
XFILLER_87_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5437__A3 _2557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7037_ clknet_leaf_12_core_clock _0298_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4249_ net2 _1736_ _1754_ _1411_ _1579_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__a221oi_4
XFILLER_247_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6398__A1 _3112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_core_clock clknet_2_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_195_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input195_A c1_sr_bus_addr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4030__C1 _1432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input362_A ic1_mem_data[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input56_A c0_o_mem_sel[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4895__A _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5428__A3 _2541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5503__B _2593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7104__CLK clknet_leaf_30_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3304__A _0896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3611__A2 _1168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output679_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7446__A net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3620_ _0871_ _1198_ _1200_ _1202_ _0874_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__a221o_1
XFILLER_174_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3551_ dmmu0.page_table\[0\]\[8\] dmmu0.page_table\[1\]\[8\] dmmu0.page_table\[2\]\[8\]
+ dmmu0.page_table\[3\]\[8\] _0897_ _0902_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__mux4_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6270_ _2801_ _3040_ vssd1 vssd1 vccd1 vccd1 _3048_ sky130_fd_sc_hd__and2_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3482_ _0879_ _1067_ _1068_ _0819_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__o31a_2
XFILLER_170_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4324__B1 _1828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5221_ net78 net77 net91 _2213_ vssd1 vssd1 vccd1 vccd1 _2426_ sky130_fd_sc_hd__or4_1
XANTENNA__4875__A1 _1989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5152_ _2249_ _2368_ _2385_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__a21o_1
XFILLER_69_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4103_ _1609_ _1610_ _1576_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__a21o_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5083_ _2332_ immu_0.page_table\[12\]\[5\] _2336_ _2343_ vssd1 vssd1 vccd1 vccd1
+ _0802_ sky130_fd_sc_hd__a31o_1
XFILLER_256_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4088__C1 _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3214__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5132__C _2373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4034_ _1423_ _1544_ _1432_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__a21o_1
XFILLER_37_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5985_ _2867_ dmmu1.page_table\[13\]\[11\] _2858_ _2874_ vssd1 vssd1 vccd1 vccd1
+ _0364_ sky130_fd_sc_hd__a31o_1
XANTENNA__6244__B _3021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5052__A1 _2316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6621__CLK clknet_leaf_53_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4936_ _2256_ vssd1 vssd1 vccd1 vccd1 _2257_ sky130_fd_sc_hd__clkbuf_4
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4867_ _1981_ _2195_ _2205_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__a21o_1
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6606_ clknet_leaf_62_core_clock _0676_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6260__A _2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3818_ net328 net382 _1360_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__mux2_2
XFILLER_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4798_ _2021_ _2155_ _2167_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__a21o_1
XFILLER_122_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6537_ clknet_leaf_44_core_clock _0607_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[14\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3749_ _1324_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_1
XFILLER_180_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6468_ _2190_ immu_1.page_table\[8\]\[5\] _3159_ vssd1 vssd1 vccd1 vccd1 _3165_ sky130_fd_sc_hd__and3_1
XFILLER_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5419_ net99 _2543_ vssd1 vssd1 vccd1 vccd1 _2548_ sky130_fd_sc_hd__and2_1
XANTENNA__7127__CLK clknet_leaf_28_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6399_ net206 _3118_ vssd1 vssd1 vccd1 vccd1 _3125_ sky130_fd_sc_hd__and2_1
XFILLER_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5604__A _2640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6419__B _3137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4618__A1 _2014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6435__A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input110_A c1_o_instr_long_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input208_A c1_sr_bus_data_o[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3794__A _0839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4402__B _1900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5514__A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4609__A1 _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6074__A3 _2922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5282__A1 _2230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6644__CLK clknet_leaf_56_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6345__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ net94 _2729_ _2745_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__a21o_1
XANTENNA__4242__C1 _1535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6794__CLK clknet_leaf_10_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4721_ _2105_ vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__buf_2
XFILLER_147_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7440_ net69 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_1
X_4652_ _2019_ _2066_ _2077_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__a21o_1
XFILLER_147_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput30 c0_o_mem_data[10] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
X_3603_ _0905_ _1180_ _1182_ net18 _1186_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__a311o_1
Xinput41 c0_o_mem_data[6] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
X_7371_ net295 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__buf_2
XFILLER_162_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4583_ _2008_ _2030_ _2035_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__a21o_1
Xinput52 c0_o_mem_high_addr[7] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
Xinput63 c0_o_req_addr[13] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_2
X_6322_ _2879_ _3079_ vssd1 vssd1 vccd1 vccd1 _3080_ sky130_fd_sc_hd__and2_1
Xinput74 c0_o_req_addr[9] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_2
X_3534_ _0869_ _1118_ _0854_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__o21a_1
Xinput85 c0_sr_bus_addr[3] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_2
Xinput96 c0_sr_bus_data_o[1] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_6
XFILLER_115_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6253_ _3036_ vssd1 vssd1 vccd1 vccd1 _3037_ sky130_fd_sc_hd__dlymetal6s2s_1
X_3465_ _0921_ _1048_ _1052_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__or3_1
XFILLER_88_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5204_ _2233_ _2409_ _2417_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__a21o_1
X_6184_ _1991_ _2982_ vssd1 vssd1 vccd1 vccd1 _2996_ sky130_fd_sc_hd__and2_1
X_3396_ dmmu0.page_table\[4\]\[3\] dmmu0.page_table\[5\]\[3\] dmmu0.page_table\[6\]\[3\]
+ dmmu0.page_table\[7\]\[3\] _0910_ _0913_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__mux4_1
XFILLER_269_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5135_ _2227_ _2369_ _2376_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__a21o_1
XFILLER_57_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5066_ _2314_ _2322_ vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__and2_1
XANTENNA__4982__B _2278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4017_ immu_1.page_table\[4\]\[2\] immu_1.page_table\[5\]\[2\] immu_1.page_table\[6\]\[2\]
+ immu_1.page_table\[7\]\[2\] _1438_ _1442_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__mux4_1
XANTENNA__6255__A _2784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5025__A1 _2301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5968_ _2805_ dmmu1.page_table\[13\]\[3\] _2859_ _2865_ vssd1 vssd1 vccd1 vccd1 _0356_
+ sky130_fd_sc_hd__a31o_1
XFILLER_12_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4919_ _1946_ vssd1 vssd1 vccd1 vccd1 _2245_ sky130_fd_sc_hd__buf_6
XFILLER_240_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5899_ _2819_ dmmu0.page_table\[6\]\[9\] _2814_ vssd1 vssd1 vccd1 vccd1 _2825_ sky130_fd_sc_hd__and3_1
XFILLER_138_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3818__S _1360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4503__A _1977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6517__CLK clknet_leaf_36_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4839__A1 _1972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input158_A c1_o_mem_long_mode vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput401 inner_wb_i_dat[6] vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_8
XFILLER_248_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5053__B _2322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6667__CLK clknet_leaf_9_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5988__B _2045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input325_A ic0_wb_cyc vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_79_core_clock clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input19_A c0_o_mem_addr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6165__A _2793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3370__S0 _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5509__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output544_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4786__C _2157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3250_ _0848_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_1
XFILLER_140_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6295__A3 _3058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4428__D_N net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6047__A3 _2902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3699__A _1280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5255__A1 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6452__B1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6940_ clknet_leaf_84_core_clock _0201_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4294__S _1408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6075__A _1897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6871_ clknet_leaf_71_core_clock _0132_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5822_ _2239_ _2767_ _2776_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__a21o_1
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5753_ _2736_ dmmu0.page_table\[4\]\[3\] _2732_ vssd1 vssd1 vccd1 vccd1 _2737_ sky130_fd_sc_hd__and3_1
XANTENNA__5419__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4704_ _2012_ _2101_ _2110_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__a21o_1
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5684_ _2235_ immu_0.high_addr_off\[5\] _2690_ vssd1 vssd1 vccd1 vccd1 _2696_ sky130_fd_sc_hd__mux2_1
XFILLER_175_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7423_ net399 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_1
X_4635_ _2067_ vssd1 vssd1 vccd1 vccd1 _2068_ sky130_fd_sc_hd__buf_2
XFILLER_190_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7354_ net308 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_2
X_4566_ _1987_ vssd1 vssd1 vccd1 vccd1 _2023_ sky130_fd_sc_hd__clkbuf_8
XFILLER_128_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6305_ _3053_ dmmu1.page_table\[4\]\[7\] _3058_ _3068_ vssd1 vssd1 vccd1 vccd1 _0490_
+ sky130_fd_sc_hd__a31o_1
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3517_ _0921_ _1098_ _1102_ _0957_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__a211o_1
X_7285_ clknet_leaf_26_core_clock _0546_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_4497_ _1939_ dmmu1.page_table\[14\]\[2\] _1964_ _1973_ vssd1 vssd1 vccd1 vccd1 _0586_
+ sky130_fd_sc_hd__a31o_1
XFILLER_277_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6236_ _2799_ _3021_ vssd1 vssd1 vccd1 vccd1 _3028_ sky130_fd_sc_hd__and2_1
XFILLER_249_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3448_ dmmu0.page_table\[6\]\[5\] dmmu0.page_table\[7\]\[5\] _0898_ vssd1 vssd1 vccd1
+ vccd1 _1036_ sky130_fd_sc_hd__mux2_1
XANTENNA__3493__A2_N _1069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4297__A2 _1799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4993__A _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _2795_ _2983_ vssd1 vssd1 vccd1 vccd1 _2987_ sky130_fd_sc_hd__and2_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ dmmu0.page_table\[4\]\[2\] dmmu0.page_table\[5\]\[2\] dmmu0.page_table\[6\]\[2\]
+ dmmu0.page_table\[7\]\[2\] _0898_ _0948_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__mux4_1
XFILLER_134_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _2363_ immu_0.page_table\[13\]\[8\] _2353_ _2364_ vssd1 vssd1 vccd1 vccd1
+ _0007_ sky130_fd_sc_hd__a31o_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ _2791_ _2944_ vssd1 vssd1 vccd1 vccd1 _2946_ sky130_fd_sc_hd__and2_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3257__A0 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5049_ _1933_ _2322_ vssd1 vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__and2_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5797__A2 _2748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5549__A2 _2623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_58_core_clock_A clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4233__A _1424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input275_A dcache_wb_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5721__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6277__A3 _3038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5485__A1 _2576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5999__A _2793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput220 dcache_mem_o_data[15] vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_4
Xinput231 dcache_wb_adr[0] vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_2
Xinput242 dcache_wb_adr[1] vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_4
XFILLER_88_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput253 dcache_wb_adr[8] vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_4
Xinput264 dcache_wb_o_dat[2] vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_6
Xinput275 dcache_wb_we vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_4
Xinput286 ic0_mem_data[18] vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_1
XFILLER_208_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5511__B _2593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput297 ic0_mem_data[28] vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4408__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3343__S0 _0891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3458__S _0896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4212__A2 _1716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7454__A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4420_ _1897_ vssd1 vssd1 vccd1 vccd1 _1910_ sky130_fd_sc_hd__buf_4
XFILLER_8_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6832__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5712__A2 _2700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput705 net705 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[9] sky130_fd_sc_hd__buf_2
XFILLER_160_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4351_ net2 _1834_ _1835_ _1854_ _1579_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__a311o_1
XFILLER_98_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3302_ net15 vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__buf_4
XFILLER_113_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7070_ clknet_leaf_4_core_clock _0331_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[6\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_4282_ immu_0.page_table\[6\]\[9\] immu_0.page_table\[7\]\[9\] _1601_ vssd1 vssd1
+ vccd1 vccd1 _1787_ sky130_fd_sc_hd__mux2_1
XFILLER_152_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_60_core_clock_A clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_6021_ _2884_ dmmu1.page_table\[12\]\[11\] _2877_ _2897_ vssd1 vssd1 vccd1 vccd1
+ _0377_ sky130_fd_sc_hd__a31o_1
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3233_ mem_dcache_arb.select net562 _0817_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__o21ai_2
XFILLER_274_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5702__A _2682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5421__B _2543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5779__A2 _2748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3222__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5140__C _2373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6440__A3 _3134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6923_ clknet_leaf_75_core_clock _0184_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6854_ clknet_leaf_70_core_clock _0115_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_5805_ _2216_ _2589_ vssd1 vssd1 vccd1 vccd1 _2766_ sky130_fd_sc_hd__nor2_1
XANTENNA__6252__B _2136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6785_ clknet_leaf_0_core_clock _0046_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[8\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3997_ immu_0.page_table\[4\]\[2\] immu_0.page_table\[5\]\[2\] immu_0.page_table\[6\]\[2\]
+ immu_0.page_table\[7\]\[2\] _1480_ _1430_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__mux4_2
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5736_ immu_1.high_addr_off\[5\] _1979_ _2720_ vssd1 vssd1 vccd1 vccd1 _2726_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_6_0_core_clock clknet_2_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_13_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5667_ _2251_ _2668_ _2685_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__a21o_1
XANTENNA__3892__A _1406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7406_ net346 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_1
X_4618_ _2014_ _2047_ _2056_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__a21o_1
XFILLER_190_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5598_ _2640_ dmmu0.page_table\[12\]\[9\] _2634_ vssd1 vssd1 vccd1 vccd1 _2645_ sky130_fd_sc_hd__and3_1
XANTENNA__5703__A2 _2700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4062__S1 _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4549_ _2010_ _2002_ _2011_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__a21o_1
XFILLER_104_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7268_ clknet_leaf_21_core_clock _0529_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6219_ _3010_ dmmu1.page_table\[7\]\[12\] _2999_ _3016_ vssd1 vssd1 vccd1 vccd1 _0456_
+ sky130_fd_sc_hd__a31o_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7199_ clknet_leaf_17_core_clock _0460_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5612__A _2640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6427__B _3137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6146__C _2962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4978__B1 _2277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6705__CLK clknet_leaf_62_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6443__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3786__B _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5059__A _1944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input392_A inner_wb_i_dat[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6855__CLK clknet_leaf_69_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input86_A c0_sr_bus_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4898__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4053__S1 _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4410__B _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3307__A _0896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5458__A1 _2562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3469__B1 _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3741__S _0847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5522__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6337__B _3079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4681__A2 _2083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5241__B _2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6422__A3 _3135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4969__B1 _2277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5630__A1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7449__A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3920_ net315 vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__inv_2
XANTENNA__5895__C _2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3696__B _1268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3851_ _1373_ net261 vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__and2_4
XFILLER_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6570_ clknet_leaf_49_core_clock _0640_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[11\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3782_ net214 _0993_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__and2_1
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5521_ _1922_ _2605_ vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__nor2_4
XFILLER_192_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3944__B2 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4601__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5452_ _2562_ immu_0.page_table\[5\]\[6\] _2557_ _2567_ vssd1 vssd1 vccd1 vccd1 _0138_
+ sky130_fd_sc_hd__a31o_1
XFILLER_145_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput502 net502 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[24] sky130_fd_sc_hd__buf_2
XANTENNA__5697__A1 _2224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4403_ _1901_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_1
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput513 net513 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[5] sky130_fd_sc_hd__buf_2
X_5383_ _2517_ immu_0.page_table\[7\]\[0\] _2525_ _2526_ vssd1 vssd1 vccd1 vccd1 _0110_
+ sky130_fd_sc_hd__a31o_1
Xoutput524 net524 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[12] sky130_fd_sc_hd__buf_2
Xoutput535 net535 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[22] sky130_fd_sc_hd__buf_2
Xoutput546 net546 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[0] sky130_fd_sc_hd__buf_2
XFILLER_172_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7122_ clknet_leaf_34_core_clock _0383_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput557 net557 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[5] sky130_fd_sc_hd__buf_2
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput568 net568 vssd1 vssd1 vccd1 vccd1 dcache_wb_err sky130_fd_sc_hd__buf_2
X_4334_ immu_0.page_table\[12\]\[10\] immu_0.page_table\[13\]\[10\] _1408_ vssd1 vssd1
+ vccd1 vccd1 _1838_ sky130_fd_sc_hd__mux2_1
XFILLER_125_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput579 net579 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[4] sky130_fd_sc_hd__buf_2
X_7053_ clknet_leaf_32_core_clock _0314_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[15\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_259_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4265_ immu_1.page_table\[6\]\[8\] immu_1.page_table\[7\]\[8\] _1453_ vssd1 vssd1
+ vccd1 vccd1 _1771_ sky130_fd_sc_hd__mux2_1
XANTENNA__7160__CLK clknet_leaf_12_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6004_ _2884_ dmmu1.page_table\[12\]\[4\] _2878_ _2887_ vssd1 vssd1 vccd1 vccd1 _0370_
+ sky130_fd_sc_hd__a31o_1
X_3216_ net228 _0824_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__and2_1
X_4196_ _1454_ _1700_ _1702_ net368 vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__o211a_1
XFILLER_227_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6728__CLK clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6413__A3 _3115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6878__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6906_ clknet_leaf_72_core_clock _0167_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6837_ clknet_leaf_68_core_clock _0098_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[9\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4188__A1 _1581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6768_ clknet_leaf_86_core_clock _0029_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5719_ _2709_ dmmu0.page_table\[2\]\[12\] _2701_ vssd1 vssd1 vccd1 vccd1 _2716_ sky130_fd_sc_hd__and3_1
XFILLER_148_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6699_ clknet_leaf_45_core_clock _0769_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5326__B _2482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input140_A c1_o_mem_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input238_A dcache_wb_adr[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5061__B _2322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6404__A3 _3116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5996__B _2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3797__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4392__S _0811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6173__A _2801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5915__A2 _2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7033__CLK clknet_leaf_13_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5517__A _1929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4421__A _1910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output457_A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4351__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5252__A _2447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4794__C _2157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4050_ immu_1.page_table\[12\]\[3\] immu_1.page_table\[13\]\[3\] _1448_ vssd1 vssd1
+ vccd1 vccd1 _1561_ sky130_fd_sc_hd__mux2_1
XANTENNA__6067__B _2924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 c0_o_instr_long_addr[1] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_4
XFILLER_36_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5603__A1 _2251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6083__A _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4952_ _2262_ immu_1.page_table\[7\]\[6\] _2259_ vssd1 vssd1 vccd1 vccd1 _2267_ sky130_fd_sc_hd__and3_1
XFILLER_205_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3500__A _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3903_ _1414_ _1415_ _1416_ vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__mux2_1
X_4883_ _2216_ vssd1 vssd1 vccd1 vccd1 _2217_ sky130_fd_sc_hd__buf_4
X_3834_ _1363_ net268 vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__and2_1
X_6622_ clknet_leaf_62_core_clock _0692_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6553_ clknet_leaf_48_core_clock _0623_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_118_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3765_ _1332_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3646__S _0847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5427__A _2310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4590__A1 _2014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5504_ _2588_ immu_0.page_table\[3\]\[5\] _2591_ _2598_ vssd1 vssd1 vccd1 vccd1 _0159_
+ sky130_fd_sc_hd__a31o_1
X_6484_ _3173_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__clkbuf_1
X_3696_ _0893_ _1268_ _1277_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__or3b_1
XANTENNA__4017__S1 _1442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5435_ _2556_ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__clkbuf_4
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5366_ _2503_ immu_0.page_table\[8\]\[4\] _2510_ _2516_ vssd1 vssd1 vccd1 vccd1 _0103_
+ sky130_fd_sc_hd__a31o_1
XFILLER_273_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4893__A2 _2219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4317_ _1496_ _1819_ _1821_ _1516_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__o211a_1
X_7105_ clknet_leaf_35_core_clock _0366_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_259_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5297_ _2249_ _2461_ _2476_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__a21o_1
XANTENNA__5162__A _2384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_274_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3528__S0 _0891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7036_ clknet_leaf_11_core_clock _0297_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4248_ _1413_ _1740_ _1744_ _1748_ _1753_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__o32a_2
XFILLER_274_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4179_ _1676_ _1682_ _1685_ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__o21a_1
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4506__A _1979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4030__B1 _1540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5373__A3 _2510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5337__A _1935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4581__A1 _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4241__A _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input188_A c1_sr_bus_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input355_A ic1_mem_data[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input49_A c0_o_mem_high_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3291__S _0865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6086__A1 _2932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4097__A0 immu_0.page_table\[8\]\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5833__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4416__A _1373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3320__A _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5946__S _2848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6010__A1 _2884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4021__B1 _1532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5364__A3 _2510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3550_ dmmu0.page_table\[4\]\[8\] dmmu0.page_table\[5\]\[8\] dmmu0.page_table\[6\]\[8\]
+ dmmu0.page_table\[7\]\[8\] _0897_ _0902_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__mux4_1
XANTENNA__6573__CLK clknet_leaf_46_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3481_ net150 dmmu1.long_off_reg\[0\] _1066_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__and3_1
XFILLER_142_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7462__A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5220_ _2253_ _2408_ _2425_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__a21o_1
XFILLER_142_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4324__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4324__B2 _1441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5151_ _2384_ dmmu0.page_table\[10\]\[10\] _2372_ vssd1 vssd1 vccd1 vccd1 _2385_
+ sky130_fd_sc_hd__and3_1
XFILLER_257_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4102_ _1576_ _1609_ _1610_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__nand3_1
X_5082_ _1940_ _2338_ vssd1 vssd1 vccd1 vccd1 _2343_ sky130_fd_sc_hd__and2_1
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3214__B _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4033_ immu_0.page_table\[0\]\[3\] immu_0.page_table\[1\]\[3\] net312 vssd1 vssd1
+ vccd1 vccd1 _1544_ sky130_fd_sc_hd__mux2_1
XFILLER_110_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7079__CLK clknet_leaf_11_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5984_ _1991_ _2860_ vssd1 vssd1 vccd1 vccd1 _2874_ sky130_fd_sc_hd__and2_1
XANTENNA__3230__A _0836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4935_ _1999_ _2255_ vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__nor2_1
XFILLER_240_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4866_ _2204_ immu_1.page_table\[3\]\[6\] _2197_ vssd1 vssd1 vccd1 vccd1 _2205_ sky130_fd_sc_hd__and3_1
XFILLER_60_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6605_ clknet_leaf_54_core_clock _0675_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6260__B _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3817_ _0812_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__buf_4
X_4797_ _2166_ immu_1.page_table\[4\]\[8\] _2157_ vssd1 vssd1 vccd1 vccd1 _2167_ sky130_fd_sc_hd__and3_1
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4699__C _2103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6536_ clknet_leaf_44_core_clock _0606_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[14\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3997__S0 _1480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3748_ net144 net39 _1322_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__mux2_2
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6467_ _1977_ _3157_ _3164_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__a21o_1
X_3679_ _0859_ _1260_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__nor2_1
XANTENNA__5107__A3 _2353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5418_ _2546_ immu_0.page_table\[6\]\[3\] _2541_ _2547_ vssd1 vssd1 vccd1 vccd1 _0124_
+ sky130_fd_sc_hd__a31o_1
X_6398_ _3112_ dmmu1.page_table\[1\]\[5\] _3116_ _3124_ vssd1 vssd1 vccd1 vccd1 _0527_
+ sky130_fd_sc_hd__a31o_1
XFILLER_217_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5349_ _2503_ immu_0.page_table\[9\]\[8\] _2495_ _2506_ vssd1 vssd1 vccd1 vccd1 _0096_
+ sky130_fd_sc_hd__a31o_1
XFILLER_101_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6068__A1 _2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4618__A2 _2047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_69_core_clock clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_275_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7019_ clknet_leaf_82_core_clock _0280_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6435__B _3137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input103_A c0_sr_bus_data_o[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6596__CLK clknet_leaf_53_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5514__B _2593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3315__A net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7221__CLK clknet_leaf_27_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4609__A2 _2047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5530__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5282__A2 _2462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6939__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4242__B1 _1747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5676__S _2690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7457__A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4720_ _2119_ vssd1 vssd1 vccd1 vccd1 _2120_ sky130_fd_sc_hd__clkbuf_4
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4793__A1 _2016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4651_ _2072_ immu_1.page_table\[11\]\[7\] _2068_ vssd1 vssd1 vccd1 vccd1 _2077_
+ sky130_fd_sc_hd__and3_1
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput20 c0_o_mem_addr[1] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
X_3602_ _0912_ _1183_ _1185_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__a21oi_1
Xinput31 c0_o_mem_data[11] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
X_4582_ _2017_ immu_1.page_table\[13\]\[2\] _2032_ vssd1 vssd1 vccd1 vccd1 _2035_
+ sky130_fd_sc_hd__and3_1
X_7370_ net294 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_2
XFILLER_174_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput42 c0_o_mem_data[7] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
Xinput53 c0_o_mem_long_mode vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_2
Xinput64 c0_o_req_addr[14] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_2
X_3533_ dmmu1.page_table\[14\]\[8\] dmmu1.page_table\[15\]\[8\] _0891_ vssd1 vssd1
+ vccd1 vccd1 _1118_ sky130_fd_sc_hd__mux2_1
X_6321_ _3078_ vssd1 vssd1 vccd1 vccd1 _3079_ sky130_fd_sc_hd__clkbuf_4
Xinput75 c0_o_req_ppl_submit vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__buf_2
Xinput86 c0_sr_bus_addr[4] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput97 c0_sr_bus_data_o[2] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__buf_4
XFILLER_143_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6252_ _2919_ _2136_ vssd1 vssd1 vccd1 vccd1 _3036_ sky130_fd_sc_hd__or2_1
X_3464_ _0909_ _1049_ _1051_ _0906_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__o211a_1
XFILLER_107_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5203_ _2416_ dmmu0.page_table\[8\]\[4\] _2411_ vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__and3_1
XFILLER_130_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6183_ _2994_ dmmu1.page_table\[8\]\[10\] _2980_ _2995_ vssd1 vssd1 vccd1 vccd1 _0441_
+ sky130_fd_sc_hd__a31o_1
X_3395_ dmmu0.page_table\[0\]\[3\] dmmu0.page_table\[1\]\[3\] dmmu0.page_table\[2\]\[3\]
+ dmmu0.page_table\[3\]\[3\] _0898_ _0913_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__mux4_1
XANTENNA__3225__A _0833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5134_ _2371_ dmmu0.page_table\[10\]\[2\] _2373_ vssd1 vssd1 vccd1 vccd1 _2376_ sky130_fd_sc_hd__and3_1
XFILLER_111_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5065_ _2300_ vssd1 vssd1 vccd1 vccd1 _2332_ sky130_fd_sc_hd__buf_4
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4016_ _1523_ _1525_ _1527_ net369 vssd1 vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__o211a_1
XFILLER_244_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6255__B _2136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5967_ _2795_ _2861_ vssd1 vssd1 vccd1 vccd1 _2865_ sky130_fd_sc_hd__and2_1
XANTENNA__3895__A _1408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4918_ _2243_ _2219_ _2244_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__a21o_1
XFILLER_279_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5898_ _1946_ _2812_ _2824_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__a21o_1
XFILLER_178_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4503__B _1970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4849_ _1999_ _2193_ vssd1 vssd1 vccd1 vccd1 _2194_ sky130_fd_sc_hd__nor2_1
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6519_ clknet_leaf_36_core_clock _0589_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7499_ net401 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__clkbuf_1
XFILLER_146_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5615__A _2655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4839__A2 _2189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5500__A3 _2591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput402 inner_wb_i_dat[7] vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_8
XFILLER_0_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5350__A _2312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4892__C _2221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6461__A1 _1967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input220_A dcache_mem_o_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input318_A ic0_wb_adr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6165__B _2983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3370__S1 _0864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6213__A1 _3010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6181__A _2931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5509__B _2593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6611__CLK clknet_leaf_53_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6356__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5260__A _2447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5255__A2 _2442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6761__CLK clknet_leaf_93_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6870_ clknet_leaf_72_core_clock _0131_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[6\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_281_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6204__A1 _2994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5821_ _2762_ dmmu0.page_table\[3\]\[6\] _2769_ vssd1 vssd1 vccd1 vccd1 _2776_ sky130_fd_sc_hd__and3_1
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7117__CLK clknet_leaf_30_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6091__A _2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4604__A _1999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5752_ _2681_ vssd1 vssd1 vccd1 vccd1 _2736_ sky130_fd_sc_hd__clkbuf_4
XFILLER_148_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4703_ _2106_ immu_1.page_table\[9\]\[4\] _2103_ vssd1 vssd1 vccd1 vccd1 _2110_ sky130_fd_sc_hd__and3_1
XFILLER_249_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3974__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5419__B _2543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5683_ _2695_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__clkbuf_1
X_7422_ net398 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_1
X_4634_ _1999_ _2064_ vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__or2_1
XANTENNA__5138__C _2373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4565_ _2021_ _2002_ _2022_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__a21o_1
X_7353_ net307 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_2
XFILLER_118_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6304_ net207 _3060_ vssd1 vssd1 vccd1 vccd1 _3068_ sky130_fd_sc_hd__and2_1
X_3516_ _0899_ _1101_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__and2_1
X_7284_ clknet_leaf_26_core_clock _0545_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4496_ _1972_ _1970_ vssd1 vssd1 vccd1 vccd1 _1973_ sky130_fd_sc_hd__and2_1
XFILLER_1_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6235_ _3026_ dmmu1.page_table\[6\]\[4\] _3019_ _3027_ vssd1 vssd1 vccd1 vccd1 _0461_
+ sky130_fd_sc_hd__a31o_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3447_ _0880_ _1026_ _1032_ _1033_ _1034_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__a32o_2
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _0899_ _0968_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__and2_1
X_6166_ _2977_ dmmu1.page_table\[8\]\[2\] _2981_ _2986_ vssd1 vssd1 vccd1 vccd1 _0433_
+ sky130_fd_sc_hd__a31o_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _2310_ _2355_ vssd1 vssd1 vccd1 vccd1 _2364_ sky130_fd_sc_hd__and2_1
XANTENNA__6266__A _2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6097_ _2932_ dmmu1.page_table\[9\]\[0\] _2942_ _2945_ vssd1 vssd1 vccd1 vccd1 _0405_
+ sky130_fd_sc_hd__a31o_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5170__A _2384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5048_ _2316_ immu_0.page_table\[14\]\[1\] _2320_ _2323_ vssd1 vssd1 vccd1 vccd1
+ _0787_ sky130_fd_sc_hd__a31o_1
XFILLER_84_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6999_ clknet_leaf_38_core_clock _0260_ vssd1 vssd1 vccd1 vccd1 immu_1.high_addr_off\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4757__A1 _2008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4514__A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5182__A1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input170_A c1_o_req_addr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input268_A dcache_wb_o_dat[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5999__B _2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput210 c1_sr_bus_we vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_1
XFILLER_248_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput221 dcache_mem_o_data[1] vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input31_A c0_o_mem_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput232 dcache_wb_adr[10] vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_2
XFILLER_209_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput243 dcache_wb_adr[20] vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_2
XFILLER_48_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4395__S _0811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput254 dcache_wb_adr[9] vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_2
XFILLER_102_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput265 dcache_wb_o_dat[3] vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__buf_6
XFILLER_236_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5080__A _1937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6434__A1 _1898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput276 ic0_mem_ack vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_1
XFILLER_236_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput287 ic0_mem_data[19] vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput298 ic0_mem_data[29] vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_1
XFILLER_90_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4408__B _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4996__A1 _1979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3343__S1 _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4460__A3 _1924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3739__S _0847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5954__S _2848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5173__A1 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput706 net706 vssd1 vssd1 vccd1 vccd1 inner_wb_sel[0] sky130_fd_sc_hd__buf_2
XANTENNA__4797__C _2157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4350_ _1844_ _1853_ _1411_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__and3b_1
XFILLER_125_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3301_ _0892_ _0893_ _0840_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__a21o_1
X_4281_ _1784_ _1785_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7470__A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6020_ _1991_ _2880_ vssd1 vssd1 vccd1 vccd1 _2897_ sky130_fd_sc_hd__and2_1
X_3232_ _0837_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_1
XFILLER_86_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3503__A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3222__B _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6922_ clknet_leaf_77_core_clock _0183_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6853_ clknet_leaf_71_core_clock _0114_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3649__S _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5804_ net95 _2747_ _2765_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__a21o_1
XANTENNA__4739__A1 _2019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6784_ clknet_leaf_89_core_clock _0045_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[8\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3996_ _1411_ _1503_ _1507_ _1479_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__a31o_1
XFILLER_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5735_ _2725_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6657__CLK clknet_leaf_42_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5666_ _2682_ dmmu0.page_table\[11\]\[11\] _2670_ vssd1 vssd1 vccd1 vccd1 _2685_
+ sky130_fd_sc_hd__and3_1
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7405_ net345 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_1
X_4617_ _2054_ immu_1.page_table\[12\]\[5\] _2049_ vssd1 vssd1 vccd1 vccd1 _2056_
+ sky130_fd_sc_hd__and3_1
XFILLER_163_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5597_ _2245_ _2632_ _2644_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__a21o_1
XFILLER_151_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4548_ _1910_ immu_1.page_table\[14\]\[3\] _2004_ vssd1 vssd1 vccd1 vccd1 _2011_
+ sky130_fd_sc_hd__and3_1
XFILLER_104_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7267_ clknet_leaf_21_core_clock _0528_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4479_ _1954_ _1957_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__or2_4
XFILLER_104_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7380__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4124__C1 _1360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6218_ _1993_ _3001_ vssd1 vssd1 vccd1 vccd1 _3016_ sky130_fd_sc_hd__and2_1
XFILLER_277_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7198_ clknet_leaf_16_core_clock _0459_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_225_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4509__A _1981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _1950_ _2959_ _2974_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__a21o_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3413__A _0855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4978__A1 _1989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6443__B _3136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4244__A _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5059__B _2322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input385_A inner_embed_mode vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input79_A c0_sr_bus_addr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5803__A _2762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3469__A1 _0957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4419__A _1909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6407__A1 _3128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4969__A1 _1967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5630__A2 _2650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3850_ _1378_ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__clkbuf_1
XFILLER_220_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3781_ _1341_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5684__S _2690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7465__A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5520_ _2603_ immu_0.page_table\[2\]\[0\] _2607_ _2608_ vssd1 vssd1 vccd1 vccd1 _0165_
+ sky130_fd_sc_hd__a31o_1
XFILLER_118_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5451_ net101 _2559_ vssd1 vssd1 vccd1 vccd1 _2567_ sky130_fd_sc_hd__and2_1
XFILLER_246_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4601__B net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4402_ _1898_ _1900_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__and2_1
Xoutput503 net503 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[25] sky130_fd_sc_hd__buf_2
XANTENNA__5697__A2 _2700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput514 net514 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[6] sky130_fd_sc_hd__buf_2
XFILLER_172_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5382_ _1926_ _2524_ vssd1 vssd1 vccd1 vccd1 _2526_ sky130_fd_sc_hd__nor2_1
Xoutput525 net525 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[13] sky130_fd_sc_hd__buf_2
Xoutput536 net536 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[23] sky130_fd_sc_hd__buf_2
Xoutput547 net547 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[10] sky130_fd_sc_hd__buf_2
XFILLER_5_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7121_ clknet_leaf_13_core_clock _0382_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput558 net558 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[6] sky130_fd_sc_hd__buf_2
X_4333_ _1478_ _1836_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__nor2_1
Xoutput569 net569 vssd1 vssd1 vccd1 vccd1 dcache_wb_i_dat[0] sky130_fd_sc_hd__buf_2
XFILLER_5_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5713__A _2709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4264_ _1763_ _1765_ _1767_ _1769_ _1553_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__o221a_2
X_7052_ clknet_leaf_32_core_clock _0313_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6110__A3 _2942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6003_ _2797_ _2881_ vssd1 vssd1 vccd1 vccd1 _2887_ sky130_fd_sc_hd__and2_1
X_3215_ _0828_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_1
X_4195_ _1446_ _1701_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__or2_1
XFILLER_39_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6905_ clknet_leaf_72_core_clock _0166_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3632__A1 _0901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6836_ clknet_leaf_69_core_clock _0097_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[9\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4999__A _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6767_ clknet_leaf_89_core_clock _0028_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3979_ _1457_ _1489_ _1491_ _1462_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__a31o_1
XFILLER_210_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5718_ _2251_ _2699_ _2715_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__a21o_1
X_6698_ clknet_leaf_45_core_clock _0768_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5137__A1 _2230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5649_ _2230_ _2669_ _2675_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__a21o_1
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5623__A _2655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6101__A3 _2942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input133_A c1_o_mem_addr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6454__A _1999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6822__CLK clknet_leaf_59_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input300_A ic0_mem_data[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3797__B _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6173__B _2983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3289__S _0865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6168__A3 _2981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5517__B _2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6340__A3 _3077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3752__S _1322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4149__A _1447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 c0_o_instr_long_addr[2] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_2
XFILLER_283_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6083__B _2924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4951_ _1979_ _2257_ _2266_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__a21o_1
XFILLER_224_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3500__B _1085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3902_ net314 vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__inv_2
XFILLER_189_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4882_ _2215_ vssd1 vssd1 vccd1 vccd1 _2216_ sky130_fd_sc_hd__buf_4
XFILLER_177_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6621_ clknet_leaf_53_core_clock _0691_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3833_ _1369_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_1
XFILLER_177_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4612__A _2038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6552_ clknet_leaf_51_core_clock _0622_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_72_core_clock_A clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3764_ net137 net32 _1322_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__mux2_4
XFILLER_192_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5427__B _2543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5503_ net100 _2593_ vssd1 vssd1 vccd1 vccd1 _2598_ sky130_fd_sc_hd__and2_1
XFILLER_185_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4590__A2 _2030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6483_ dmmu1.long_off_reg\[0\] _1995_ _3172_ vssd1 vssd1 vccd1 vccd1 _3173_ sky130_fd_sc_hd__mux2_1
XFILLER_145_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3695_ _0872_ _1270_ _1272_ _1276_ net123 vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__a311o_2
XFILLER_257_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3228__A _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5146__C _2373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5434_ _1929_ _2555_ vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__or2_1
XFILLER_279_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6331__A3 _3077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5365_ _1937_ _2512_ vssd1 vssd1 vccd1 vccd1 _2516_ sky130_fd_sc_hd__and2_1
XFILLER_259_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3662__S _1169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5443__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7104_ clknet_leaf_30_core_clock _0365_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[13\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_4316_ _1584_ _1820_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__or2_1
XFILLER_141_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5296_ _2473_ dmmu0.page_table\[14\]\[10\] _2463_ vssd1 vssd1 vccd1 vccd1 _2476_
+ sky130_fd_sc_hd__and3_1
XFILLER_275_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_59_core_clock clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_core_clock
+ sky130_fd_sc_hd__clkbuf_16
X_7035_ clknet_leaf_12_core_clock _0296_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3528__S1 _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4247_ _1479_ _1750_ _1752_ _1434_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__a31o_1
XANTENNA__4059__A inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6845__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4178_ _1683_ _1684_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__nand2_1
XFILLER_262_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3898__A _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_255_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6274__A _2891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6398__A3 _3116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4506__B _1970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6995__CLK clknet_leaf_1_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6819_ clknet_leaf_68_core_clock _0080_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4030__A1 _1424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5337__B _2497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4581__A2 _2030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3572__S _1146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input250_A dcache_wb_adr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input348_A ic1_mem_data[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4097__A1 immu_0.page_table\[9\]\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6184__A _1991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5597__A1 _2245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7000__CLK clknet_leaf_37_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4416__B net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5349__A1 _2503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7150__CLK clknet_leaf_35_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5528__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4432__A _1921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4021__A1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6718__CLK clknet_leaf_62_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4309__C1 _1516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3480_ net150 dmmu1.long_off_reg\[0\] _1066_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__a21oi_1
XFILLER_155_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6359__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5150_ _2370_ vssd1 vssd1 vccd1 vccd1 _2384_ sky130_fd_sc_hd__buf_2
XFILLER_269_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4101_ net6 immu_0.high_addr_off\[1\] vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__or2_1
XFILLER_243_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5081_ _2332_ immu_0.page_table\[12\]\[4\] _2336_ _2342_ vssd1 vssd1 vccd1 vccd1
+ _0801_ sky130_fd_sc_hd__a31o_1
XFILLER_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4088__A1 _1462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4032_ immu_0.page_table\[2\]\[3\] immu_0.page_table\[3\]\[3\] _1472_ vssd1 vssd1
+ vccd1 vccd1 _1543_ sky130_fd_sc_hd__mux2_1
XFILLER_244_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6094__A _1968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5588__A1 _2233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5983_ _2867_ dmmu1.page_table\[13\]\[10\] _2858_ _2873_ vssd1 vssd1 vccd1 vccd1
+ _0363_ sky130_fd_sc_hd__a31o_1
XFILLER_252_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5052__A3 _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4934_ _2063_ _2117_ vssd1 vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__or2_2
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4865_ _2105_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__buf_4
XFILLER_268_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3657__S _0896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5438__A _1922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6604_ clknet_leaf_53_core_clock _0674_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3816_ _1359_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4342__A _1424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4796_ _2105_ vssd1 vssd1 vccd1 vccd1 _2166_ sky130_fd_sc_hd__buf_2
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6535_ clknet_leaf_45_core_clock _0605_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[14\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3747_ _1323_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5760__A1 _2239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3997__S1 _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6466_ _2971_ immu_1.page_table\[8\]\[4\] _3159_ vssd1 vssd1 vccd1 vccd1 _3164_ sky130_fd_sc_hd__and3_1
X_3678_ dmmu1.page_table\[8\]\[11\] dmmu1.page_table\[9\]\[11\] _1146_ vssd1 vssd1
+ vccd1 vccd1 _1260_ sky130_fd_sc_hd__mux2_1
XFILLER_118_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5417_ net98 _2543_ vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__and2_1
XANTENNA__5512__A1 _2588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6397_ net205 _3118_ vssd1 vssd1 vccd1 vccd1 _3124_ sky130_fd_sc_hd__and2_1
XFILLER_217_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5348_ _2310_ _2497_ vssd1 vssd1 vccd1 vccd1 _2506_ sky130_fd_sc_hd__and2_1
XFILLER_87_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5279_ _2458_ dmmu0.page_table\[14\]\[2\] _2464_ vssd1 vssd1 vccd1 vccd1 _2467_ sky130_fd_sc_hd__and3_1
XANTENNA__5901__A _2819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7018_ clknet_leaf_4_core_clock _0279_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[4\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__7023__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4517__A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7173__CLK clknet_leaf_12_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3567__S _1146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5348__A _2310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4252__A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input298_A ic0_mem_data[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5751__A1 _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3762__A0 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input61_A c0_o_req_addr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6179__A _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5811__A _2762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_0_0_core_clock clknet_1_0_1_core_clock vssd1 vssd1 vccd1 vccd1 clknet_2_0_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_253_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4242__A1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4793__A2 _2155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6361__B _3098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3477__S _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5258__A _2447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4162__A _1447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4650_ _2016_ _2066_ _2076_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__a21o_1
XFILLER_174_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 c0_o_instr_long_addr[5] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_2
X_3601_ _0908_ _1184_ _0905_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__a21o_1
Xinput21 c0_o_mem_addr[2] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
X_4581_ _2006_ _2030_ _2034_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__a21o_1
Xinput32 c0_o_mem_data[12] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 c0_o_mem_data[8] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
Xinput54 c0_o_mem_req vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XANTENNA__6690__CLK clknet_leaf_58_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7473__A net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6320_ _2784_ _2193_ vssd1 vssd1 vccd1 vccd1 _3078_ sky130_fd_sc_hd__nor2_1
XFILLER_143_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3532_ _0863_ _1116_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__or2_1
Xinput65 c0_o_req_addr[15] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__buf_2
Xinput76 c0_sr_bus_addr[0] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_2
XFILLER_155_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput87 c0_sr_bus_addr[5] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
Xinput98 c0_sr_bus_data_o[3] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_4
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6251_ _3026_ dmmu1.page_table\[6\]\[12\] _3018_ _3035_ vssd1 vssd1 vccd1 vccd1 _0469_
+ sky130_fd_sc_hd__a31o_1
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6089__A _1993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3463_ _0913_ _1050_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__or2_1
XFILLER_88_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5202_ _2370_ vssd1 vssd1 vccd1 vccd1 _2416_ sky130_fd_sc_hd__clkbuf_4
X_6182_ _2895_ _2982_ vssd1 vssd1 vccd1 vccd1 _2995_ sky130_fd_sc_hd__and2_1
XFILLER_276_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7046__CLK clknet_leaf_32_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3394_ _0874_ _0880_ _0983_ _0840_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__a31o_2
XFILLER_257_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5133_ _2224_ _2369_ _2375_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__a21o_1
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5064_ _2316_ immu_0.page_table\[14\]\[9\] _2320_ _2331_ vssd1 vssd1 vccd1 vccd1
+ _0795_ sky130_fd_sc_hd__a31o_1
XFILLER_229_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4015_ _1442_ _1526_ vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__or2_1
XFILLER_37_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4337__A _1570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5025__A3 _2298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5966_ _2805_ dmmu1.page_table\[13\]\[2\] _2859_ _2864_ vssd1 vssd1 vccd1 vccd1 _0355_
+ sky130_fd_sc_hd__a31o_1
XFILLER_240_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4917_ _2237_ dmmu0.page_table\[0\]\[7\] _2221_ vssd1 vssd1 vccd1 vccd1 _2244_ sky130_fd_sc_hd__and3_1
XANTENNA__5981__A1 _2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5897_ _2819_ dmmu0.page_table\[6\]\[8\] _2814_ vssd1 vssd1 vccd1 vccd1 _2824_ sky130_fd_sc_hd__and3_1
XANTENNA__5168__A _2384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4848_ net190 net189 _2063_ vssd1 vssd1 vccd1 vccd1 _2193_ sky130_fd_sc_hd__or3_4
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4779_ _2156_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__buf_2
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6518_ clknet_leaf_43_core_clock _0588_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7498_ net400 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6449_ mem_dcache_arb.transfer_active vssd1 vssd1 vccd1 vccd1 _3153_ sky130_fd_sc_hd__inv_2
XFILLER_164_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput403 inner_wb_i_dat[8] vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_8
XFILLER_87_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5631__A _2655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5350__B _2497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6461__A2 _3157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4472__A1 _1939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6563__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input213_A dcache_mem_exception vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6462__A _2971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5078__A _1935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4083__S0 _1439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7069__CLK clknet_leaf_4_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output432_A net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3760__S _1322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5541__A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6356__B _3098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4157__A _1581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4463__A1 _1939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7468__A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5820_ _2235_ _2767_ _2775_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__a21o_1
XFILLER_234_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5751_ _2226_ _2730_ _2735_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__a21o_1
XANTENNA__6091__B _2099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4604__B _2045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_core_clock_A clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_222_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4702_ _2010_ _2101_ _2109_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__a21o_1
X_5682_ _2232_ immu_0.high_addr_off\[4\] _2690_ vssd1 vssd1 vccd1 vccd1 _2695_ sky130_fd_sc_hd__mux2_1
XFILLER_30_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7421_ net397 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_1
XFILLER_175_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4633_ _2065_ vssd1 vssd1 vccd1 vccd1 _2066_ sky130_fd_sc_hd__clkbuf_4
XFILLER_147_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3935__S _1448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7352_ net306 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_2
XFILLER_118_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4564_ _2017_ immu_1.page_table\[14\]\[8\] _2004_ vssd1 vssd1 vccd1 vccd1 _2022_
+ sky130_fd_sc_hd__and3_1
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6303_ _3053_ dmmu1.page_table\[4\]\[6\] _3058_ _3067_ vssd1 vssd1 vccd1 vccd1 _0489_
+ sky130_fd_sc_hd__a31o_1
X_3515_ _1099_ _1100_ _0917_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__mux2_1
X_7283_ clknet_leaf_25_core_clock _0544_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4495_ net202 vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__buf_6
X_6234_ _2797_ _3021_ vssd1 vssd1 vccd1 vccd1 _3027_ sky130_fd_sc_hd__and2_1
XANTENNA__6140__A1 _2239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3446_ net158 _0878_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__and2_2
XFILLER_170_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _2793_ _2983_ vssd1 vssd1 vccd1 vccd1 _2986_ sky130_fd_sc_hd__and2_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ dmmu0.page_table\[12\]\[2\] dmmu0.page_table\[13\]\[2\] dmmu0.page_table\[14\]\[2\]
+ dmmu0.page_table\[15\]\[2\] _0898_ _0948_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__mux4_1
XANTENNA__4993__C _2282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _2300_ vssd1 vssd1 vccd1 vccd1 _2363_ sky130_fd_sc_hd__buf_4
XANTENNA__6586__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6266__B _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6096_ _2879_ _2944_ vssd1 vssd1 vccd1 vccd1 _2945_ sky130_fd_sc_hd__and2_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5047_ _1928_ _2322_ vssd1 vssd1 vccd1 vccd1 _2323_ sky130_fd_sc_hd__and2_1
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7378__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6998_ clknet_leaf_39_core_clock _0259_ vssd1 vssd1 vccd1 vccd1 immu_1.high_addr_off\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5949_ _2853_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5954__A1 _1944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4757__A2 _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4065__S0 _1479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4530__A _1995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5182__A2 _2390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input163_A c1_o_req_active vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5485__A3 _2574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput200 c1_sr_bus_data_o[12] vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_2
XFILLER_88_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput211 core_reset vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_6
XANTENNA__5361__A _1933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput222 dcache_mem_o_data[2] vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_4
XFILLER_248_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput233 dcache_wb_adr[11] vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_2
XFILLER_76_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_core_clock_A core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input330_A ic1_mem_ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput244 dcache_wb_adr[21] vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_2
Xinput255 dcache_wb_cyc vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__buf_4
Xinput266 dcache_wb_o_dat[4] vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_6
XANTENNA__5080__B _2338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput277 ic0_mem_data[0] vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input24_A c0_o_mem_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput288 ic0_mem_data[1] vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_1
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput299 ic0_mem_data[2] vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4408__C net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4996__A2 _2280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4705__A _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6198__A1 _2994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_2_core_clock_A clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5536__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4440__A _1921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_77_core_clock_A clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_144_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6370__A1 _3101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5173__A2 _2390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput707 net707 vssd1 vssd1 vccd1 vccd1 inner_wb_sel[1] sky130_fd_sc_hd__buf_2
XFILLER_144_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3300_ net106 net158 _0879_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__o21ai_2
XANTENNA__6122__A1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4280_ _1733_ _1735_ _1732_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__o21bai_1
XFILLER_152_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3231_ net220 _0835_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__and2_2
XANTENNA__6367__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5271__A _2217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5702__C _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6921_ clknet_leaf_57_core_clock _0182_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_282_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4615__A _2054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6852_ clknet_leaf_68_core_clock _0113_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7234__CLK clknet_leaf_26_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5803_ _2762_ dmmu0.page_table\[13\]\[12\] _2750_ vssd1 vssd1 vccd1 vccd1 _2765_
+ sky130_fd_sc_hd__and3_1
XFILLER_250_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6783_ clknet_leaf_90_core_clock _0044_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[8\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5936__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4739__A2 _2120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3995_ _1420_ _1504_ _1506_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__a21o_1
XFILLER_250_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5734_ immu_1.high_addr_off\[4\] _1977_ _2720_ vssd1 vssd1 vccd1 vccd1 _2725_ sky130_fd_sc_hd__mux2_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5665_ _2249_ _2668_ _2684_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__a21o_1
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7404_ net344 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_1
X_4616_ _2012_ _2047_ _2055_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__a21o_1
XFILLER_190_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5596_ _2640_ dmmu0.page_table\[12\]\[8\] _2634_ vssd1 vssd1 vccd1 vccd1 _2644_ sky130_fd_sc_hd__and3_1
X_4547_ _1974_ vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__buf_6
XFILLER_190_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7266_ clknet_leaf_20_core_clock _0527_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4478_ net710 _1956_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__or2_1
XFILLER_143_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6217_ _3010_ dmmu1.page_table\[7\]\[11\] _2999_ _3015_ vssd1 vssd1 vccd1 vccd1 _0455_
+ sky130_fd_sc_hd__a31o_1
XFILLER_104_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3429_ _1012_ _1014_ _1017_ _0921_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__a22o_1
XFILLER_77_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7197_ clknet_leaf_28_core_clock _0458_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4675__A1 _2012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5181__A _2400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5612__C _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6148_ _2971_ dmmu0.page_table\[1\]\[10\] _2961_ vssd1 vssd1 vccd1 vccd1 _2974_ sky130_fd_sc_hd__and3_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4509__B _1970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6079_ _2803_ _2924_ vssd1 vssd1 vccd1 vccd1 _2934_ sky130_fd_sc_hd__and2_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4006__B_N _1448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5927__A1 _2242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6601__CLK clknet_leaf_54_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3938__B1 _1451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0_0_core_clock_A clknet_1_0_1_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3402__A2 _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3575__S _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5356__A _1926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input280_A ic0_mem_data[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input378_A ic1_wb_adr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6104__A1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4115__B1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5458__A3 _2557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7107__CLK clknet_leaf_36_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4666__A1 _1996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5091__A _2312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7257__CLK clknet_leaf_25_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4969__A2 _2274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4435__A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3780_ net212 _0993_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__and2_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3485__S _0918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5266__A _2370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5450_ _2562_ immu_0.page_table\[5\]\[5\] _2557_ _2566_ vssd1 vssd1 vccd1 vccd1 _0137_
+ sky130_fd_sc_hd__a31o_1
XFILLER_157_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4401_ net255 _1899_ _0811_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__mux2_4
XFILLER_172_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput504 net504 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[26] sky130_fd_sc_hd__buf_2
XFILLER_145_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5381_ _2524_ vssd1 vssd1 vccd1 vccd1 _2525_ sky130_fd_sc_hd__clkbuf_4
Xoutput515 net515 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[7] sky130_fd_sc_hd__buf_2
Xoutput526 net526 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[14] sky130_fd_sc_hd__buf_2
Xoutput537 net537 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[2] sky130_fd_sc_hd__buf_2
XFILLER_160_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7120_ clknet_leaf_14_core_clock _0381_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput548 net548 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[11] sky130_fd_sc_hd__buf_2
X_4332_ immu_0.page_table\[14\]\[10\] immu_0.page_table\[15\]\[10\] _1480_ vssd1 vssd1
+ vccd1 vccd1 _1836_ sky130_fd_sc_hd__mux2_1
XFILLER_113_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput559 net559 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[7] sky130_fd_sc_hd__buf_2
XFILLER_5_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7051_ clknet_leaf_36_core_clock _0312_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_49_core_clock clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_core_clock
+ sky130_fd_sc_hd__clkbuf_16
X_4263_ _1581_ _1768_ _1516_ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__o21ai_1
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6002_ _2884_ dmmu1.page_table\[12\]\[3\] _2878_ _2886_ vssd1 vssd1 vccd1 vccd1 _0369_
+ sky130_fd_sc_hd__a31o_1
XFILLER_274_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3214_ net227 _0824_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__and2_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4194_ immu_1.page_table\[14\]\[7\] immu_1.page_table\[15\]\[7\] net366 vssd1 vssd1
+ vccd1 vccd1 _1701_ sky130_fd_sc_hd__mux2_1
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6624__CLK clknet_leaf_54_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6904_ clknet_leaf_79_core_clock _0165_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6835_ clknet_leaf_69_core_clock _0096_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[9\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6766_ clknet_leaf_87_core_clock _0027_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3978_ _1447_ net368 _1490_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__or3_1
XFILLER_138_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5717_ _2709_ dmmu0.page_table\[2\]\[11\] _2701_ vssd1 vssd1 vccd1 vccd1 _2715_ sky130_fd_sc_hd__and3_1
X_6697_ clknet_leaf_42_core_clock _0767_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5176__A _2370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4080__A _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6334__A1 _3085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5137__A2 _2369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5648_ _2666_ dmmu0.page_table\[11\]\[3\] _2671_ vssd1 vssd1 vccd1 vccd1 _2675_ sky130_fd_sc_hd__and3_1
XFILLER_163_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_88_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5579_ _2473_ dmmu0.page_table\[12\]\[0\] _2634_ vssd1 vssd1 vccd1 vccd1 _2635_ sky130_fd_sc_hd__and3_1
XANTENNA__7391__A net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7249_ clknet_leaf_24_core_clock _0510_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4648__A1 _2014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input126_A c1_o_mem_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6470__A _2190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input91_A c0_sr_bus_addr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5086__A _1944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6325__A1 _3069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4639__A1 _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3334__A net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5252__C _2445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6647__CLK clknet_leaf_43_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 c0_o_instr_long_addr[3] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_2
XFILLER_264_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5064__A1 _2316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4950_ _2262_ immu_1.page_table\[7\]\[5\] _2259_ vssd1 vssd1 vccd1 vccd1 _2266_ sky130_fd_sc_hd__and3_1
XANTENNA__4165__A _1441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4272__C1 _1451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4811__A1 _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3901_ immu_0.page_table\[0\]\[0\] immu_0.page_table\[1\]\[0\] immu_0.page_table\[2\]\[0\]
+ immu_0.page_table\[3\]\[0\] _1407_ net313 vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__mux4_1
XANTENNA__6797__CLK clknet_leaf_10_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4881_ _1920_ _2214_ vssd1 vssd1 vccd1 vccd1 _2215_ sky130_fd_sc_hd__or2_2
XFILLER_220_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6620_ clknet_leaf_53_core_clock _0690_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3832_ _1363_ net267 vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__and2_1
XANTENNA__6380__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6551_ clknet_leaf_51_core_clock _0621_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3763_ _1331_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_2
XFILLER_158_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5502_ _2588_ immu_0.page_table\[3\]\[4\] _2591_ _2597_ vssd1 vssd1 vccd1 vccd1 _0158_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__6316__A1 _3069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6482_ _1954_ _2719_ vssd1 vssd1 vccd1 vccd1 _3172_ sky130_fd_sc_hd__nor2_8
XFILLER_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3694_ _0868_ _1273_ _1275_ _0854_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__o211a_1
XFILLER_145_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5433_ _2350_ _2439_ vssd1 vssd1 vccd1 vccd1 _2555_ sky130_fd_sc_hd__or2_4
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5724__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5364_ _2503_ immu_0.page_table\[8\]\[3\] _2510_ _2515_ vssd1 vssd1 vccd1 vccd1 _0102_
+ sky130_fd_sc_hd__a31o_1
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7103_ clknet_leaf_30_core_clock _0364_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[13\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_273_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4315_ immu_1.page_table\[6\]\[9\] immu_1.page_table\[7\]\[9\] _1493_ vssd1 vssd1
+ vccd1 vccd1 _1820_ sky130_fd_sc_hd__mux2_1
XANTENNA__5443__B _2559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5295_ _2247_ _2462_ _2475_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__a21o_1
XFILLER_87_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5162__C _2392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7034_ clknet_leaf_13_core_clock _0295_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_247_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4246_ _1478_ _1751_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__or2_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4177_ net113 immu_1.high_addr_off\[3\] vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__or2_1
XFILLER_255_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3898__B _1411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6274__B _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4802__A1 _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7386__A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout710_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6290__A _2879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4803__A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6818_ clknet_leaf_59_core_clock _0079_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6749_ clknet_leaf_87_core_clock _0010_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4014__S _1448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4869__A1 _1983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input243_A dcache_wb_adr[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6184__B _2982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5597__A2 _2632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5809__A _2762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4713__A _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6010__A3 _2878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_core_clock_A clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_174_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4021__A2 _1508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5544__A _1921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6359__B _3098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4100_ net6 immu_0.high_addr_off\[1\] vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__nand2_1
X_5080_ _1937_ _2338_ vssd1 vssd1 vccd1 vccd1 _2342_ sky130_fd_sc_hd__and2_1
XFILLER_256_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4088__A2 _1588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4031_ _1413_ _1410_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__nand2_1
XANTENNA__6375__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3391__S0 _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6094__B _2099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5982_ _1989_ _2860_ vssd1 vssd1 vccd1 vccd1 _2873_ sky130_fd_sc_hd__and2_1
XANTENNA__5588__A2 _2632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3599__A1 dmmu0.page_table\[3\]\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4933_ _2253_ _2218_ _2254_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__a21o_1
XFILLER_178_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5719__A _2709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4623__A _2054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4864_ _1979_ _2195_ _2203_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__a21o_1
X_6603_ clknet_leaf_41_core_clock _0673_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[6\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3815_ net213 _0840_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__and2_1
XANTENNA__5438__B _2555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4795_ _2019_ _2155_ _2165_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__a21o_1
XFILLER_165_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3239__A _0842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6534_ clknet_leaf_47_core_clock _0604_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3746_ net143 net38 _1322_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__mux2_1
XFILLER_118_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5760__A2 _2730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6465_ _1974_ _3157_ _3163_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__a21o_1
X_3677_ _1256_ _1257_ _1255_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__a21oi_1
XFILLER_133_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5416_ _2300_ vssd1 vssd1 vccd1 vccd1 _2546_ sky130_fd_sc_hd__clkbuf_4
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6396_ _3112_ dmmu1.page_table\[1\]\[4\] _3116_ _3123_ vssd1 vssd1 vccd1 vccd1 _0526_
+ sky130_fd_sc_hd__a31o_1
X_5347_ _2503_ immu_0.page_table\[9\]\[7\] _2495_ _2505_ vssd1 vssd1 vccd1 vccd1 _0095_
+ sky130_fd_sc_hd__a31o_1
XFILLER_102_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6068__A3 _2922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5278_ _2224_ _2462_ _2466_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__a21o_1
XANTENNA__5276__A1 _2211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7017_ clknet_leaf_17_core_clock _0278_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[4\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_247_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4229_ _1708_ _1709_ _1707_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__a21boi_2
XANTENNA__6285__A _2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3382__S0 _0898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5629__A _2655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4533__A _1998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5348__B _2497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_core_clock_A clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_129_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinterconnect_inner_730 vssd1 vssd1 vccd1 vccd1 interconnect_inner_730/HI c1_i_core_int_sreg[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4003__A2 _1509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input193_A c1_sr_bus_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5751__A2 _2730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input360_A ic1_mem_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6179__B _2983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input54_A c0_o_mem_req vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5811__B dmmu0.page_table\[3\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6195__A _2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3373__S0 _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5019__A1 _2301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3758__S _1322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4242__A2 _1745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5539__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4443__A _1928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output677_A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6835__CLK clknet_leaf_69_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3600_ dmmu0.page_table\[0\]\[9\] dmmu0.page_table\[1\]\[9\] _0895_ vssd1 vssd1 vccd1
+ vccd1 _1184_ sky130_fd_sc_hd__mux2_1
Xinput11 c0_o_instr_long_addr[6] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_2
X_4580_ _2017_ immu_1.page_table\[13\]\[1\] _2032_ vssd1 vssd1 vccd1 vccd1 _2034_
+ sky130_fd_sc_hd__and3_1
Xinput22 c0_o_mem_addr[3] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput33 c0_o_mem_data[13] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
Xinput44 c0_o_mem_data[9] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3531_ dmmu1.page_table\[12\]\[8\] dmmu1.page_table\[13\]\[8\] _0857_ vssd1 vssd1
+ vccd1 vccd1 _1116_ sky130_fd_sc_hd__mux2_1
Xinput55 c0_o_mem_sel[0] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput66 c0_o_req_addr[1] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__buf_2
Xinput77 c0_sr_bus_addr[10] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput88 c0_sr_bus_addr[6] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_1
XFILLER_155_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6250_ _1993_ _3020_ vssd1 vssd1 vccd1 vccd1 _3035_ sky130_fd_sc_hd__and2_1
Xinput99 c0_sr_bus_data_o[4] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3462_ dmmu0.page_table\[12\]\[5\] dmmu0.page_table\[13\]\[5\] _0900_ vssd1 vssd1
+ vccd1 vccd1 _1050_ sky130_fd_sc_hd__mux2_1
XFILLER_254_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5201_ _2230_ _2409_ _2415_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__a21o_1
XANTENNA__6985__CLK clknet_leaf_7_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6181_ _2931_ vssd1 vssd1 vccd1 vccd1 _2994_ sky130_fd_sc_hd__buf_4
X_3393_ _0981_ _0982_ _0855_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__mux2_1
XFILLER_269_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5132_ _2371_ dmmu0.page_table\[10\]\[1\] _2373_ vssd1 vssd1 vccd1 vccd1 _2375_ sky130_fd_sc_hd__and3_1
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5063_ _2312_ _2322_ vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__and2_1
XFILLER_257_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4014_ immu_1.page_table\[12\]\[2\] immu_1.page_table\[13\]\[2\] _1448_ vssd1 vssd1
+ vccd1 vccd1 _1526_ sky130_fd_sc_hd__mux2_1
XFILLER_265_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_84_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_65_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5965_ _2793_ _2861_ vssd1 vssd1 vccd1 vccd1 _2864_ sky130_fd_sc_hd__and2_1
XANTENNA__5430__A1 _2546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5449__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4353__A _1523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4916_ _2242_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__buf_4
X_5896_ _2242_ _2812_ _2823_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__a21o_1
XFILLER_178_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4847_ _1989_ _2188_ _2191_ immu_1.page_table\[1\]\[10\] vssd1 vssd1 vccd1 vccd1
+ _0717_ sky130_fd_sc_hd__o22a_1
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4778_ _2084_ _2153_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__or2_1
XFILLER_119_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3729_ dmmu1.page_table\[8\]\[12\] dmmu1.page_table\[9\]\[12\] dmmu1.page_table\[10\]\[12\]
+ dmmu1.page_table\[11\]\[12\] _1146_ _0859_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__mux4_1
X_6517_ clknet_leaf_36_core_clock _0587_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7497_ net399 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_1
XFILLER_106_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5615__C _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6448_ net211 _0810_ _0819_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__nor3_1
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6379_ _1910_ vssd1 vssd1 vccd1 vccd1 _3112_ sky130_fd_sc_hd__clkbuf_4
Xinput404 inner_wb_i_dat[9] vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_8
XANTENNA__5249__A1 _2227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7140__CLK clknet_leaf_29_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6213__A3 _3000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input206_A c1_sr_bus_data_o[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7290__CLK clknet_leaf_92_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5359__A _1928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6858__CLK clknet_leaf_69_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5078__B _2338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4083__S1 _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5260__C _2445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6452__A3 _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6204__A3 _3000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3488__S _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5269__A _2458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5750_ _2709_ dmmu0.page_table\[4\]\[2\] _2732_ vssd1 vssd1 vccd1 vccd1 _2735_ sky130_fd_sc_hd__and3_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4701_ _2106_ immu_1.page_table\[9\]\[3\] _2103_ vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__and3_1
XFILLER_249_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3974__A1 _1451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5681_ _2694_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__clkbuf_1
X_4632_ _2000_ _2064_ vssd1 vssd1 vccd1 vccd1 _2065_ sky130_fd_sc_hd__nor2_1
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7420_ net396 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_1
XANTENNA__7013__CLK clknet_leaf_37_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3726__A1 _0869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4563_ _1985_ vssd1 vssd1 vccd1 vccd1 _2021_ sky130_fd_sc_hd__buf_4
X_7351_ net305 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_2
XFILLER_116_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4112__S _1493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6302_ net206 _3060_ vssd1 vssd1 vccd1 vccd1 _3067_ sky130_fd_sc_hd__and2_1
X_3514_ dmmu0.page_table\[8\]\[7\] dmmu0.page_table\[9\]\[7\] dmmu0.page_table\[10\]\[7\]
+ dmmu0.page_table\[11\]\[7\] _0896_ _0901_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__mux4_1
XFILLER_155_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7282_ clknet_leaf_24_core_clock _0543_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4494_ _1939_ dmmu1.page_table\[14\]\[1\] _1964_ _1971_ vssd1 vssd1 vccd1 vccd1 _0585_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__5479__A1 _2576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6233_ _2931_ vssd1 vssd1 vccd1 vccd1 _3026_ sky130_fd_sc_hd__buf_4
XFILLER_143_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3445_ net150 dmmu1.long_off_reg\[0\] vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__xor2_1
XANTENNA__6140__A2 _2960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7163__CLK clknet_leaf_9_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6164_ _2977_ dmmu1.page_table\[8\]\[1\] _2981_ _2985_ vssd1 vssd1 vccd1 vccd1 _0432_
+ sky130_fd_sc_hd__a31o_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3376_ _0881_ _0880_ _0966_ _0840_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__a31o_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__B _2559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5115_ _2347_ immu_0.page_table\[13\]\[7\] _2353_ _2362_ vssd1 vssd1 vccd1 vccd1
+ _0006_ sky130_fd_sc_hd__a31o_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _2943_ vssd1 vssd1 vccd1 vccd1 _2944_ sky130_fd_sc_hd__clkbuf_4
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3252__A _0849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5170__C _2392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5046_ _1930_ _2318_ vssd1 vssd1 vccd1 vccd1 _2322_ sky130_fd_sc_hd__nor2_4
XFILLER_245_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5651__A1 _2233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5403__A1 _2531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6997_ clknet_leaf_62_core_clock _0258_ vssd1 vssd1 vccd1 vccd1 icache_arbiter.o_sel_sig
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5179__A _2400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5948_ dmmu0.long_off_reg\[4\] _1937_ _2848_ vssd1 vssd1 vccd1 vccd1 _2853_ sky130_fd_sc_hd__mux2_1
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5879_ _2813_ vssd1 vssd1 vccd1 vccd1 _2814_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__7394__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5907__A _2216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4022__S _0811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3861__S _1360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5642__A _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input156_A c1_o_mem_high_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6530__CLK clknet_leaf_42_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput201 c1_sr_bus_data_o[1] vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_4
XFILLER_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3350__C1 _0855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5361__B _2512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput212 dcache_mem_ack vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_2
XANTENNA__5890__A1 _2232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput223 dcache_mem_o_data[3] vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput234 dcache_wb_adr[12] vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_2
XFILLER_75_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput245 dcache_wb_adr[22] vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_4
XFILLER_248_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput256 dcache_wb_o_dat[0] vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_6
XFILLER_124_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput267 dcache_wb_o_dat[5] vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_6
XANTENNA_input323_A ic0_wb_adr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6434__A3 _3135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput278 ic0_mem_data[10] vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput289 ic0_mem_data[20] vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_1
XFILLER_263_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input17_A c0_o_mem_addr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6680__CLK clknet_leaf_54_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7036__CLK clknet_leaf_11_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5817__A _2762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4721__A _2105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput708 net708 vssd1 vssd1 vccd1 vccd1 inner_wb_stb sky130_fd_sc_hd__buf_2
XANTENNA_output542_A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_39_core_clock clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_152_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3230_ _0836_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4133__A1 _1535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6367__B _3098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5271__B _2318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5881__A1 _2210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4168__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6920_ clknet_leaf_76_core_clock _0181_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_254_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3927__A_N net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6851_ clknet_leaf_69_core_clock _0112_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_207_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5802_ net94 _2747_ _2764_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__a21o_1
XFILLER_222_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6782_ clknet_leaf_89_core_clock _0043_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3994_ _1424_ _1505_ _1434_ vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__a21o_1
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3947__A1 _1460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5733_ _2724_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5664_ _2682_ dmmu0.page_table\[11\]\[10\] _2670_ vssd1 vssd1 vccd1 vccd1 _2684_
+ sky130_fd_sc_hd__and3_1
XFILLER_129_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_78_core_clock clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_core_clock
+ sky130_fd_sc_hd__clkbuf_16
X_7403_ net343 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_1
XFILLER_175_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4615_ _2054_ immu_1.page_table\[12\]\[4\] _2049_ vssd1 vssd1 vccd1 vccd1 _2055_
+ sky130_fd_sc_hd__and3_1
XFILLER_163_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5595_ _2243_ _2632_ _2643_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__a21o_1
XFILLER_209_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3247__A _0846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4546_ _2008_ _2002_ _2009_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__a21o_1
XANTENNA__6553__CLK clknet_leaf_48_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7265_ clknet_leaf_24_core_clock _0526_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4477_ net191 _1955_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__or2_1
XFILLER_1_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5462__A _1929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6216_ _1991_ _3001_ vssd1 vssd1 vccd1 vccd1 _3015_ sky130_fd_sc_hd__and2_1
X_3428_ _1015_ _1016_ _0906_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__mux2_1
XFILLER_131_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7196_ clknet_leaf_16_core_clock _0457_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_277_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4675__A2 _2083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A c0_o_instr_long_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6147_ _1948_ _2960_ _2973_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__a21o_1
X_3359_ dmmu0.page_table\[2\]\[1\] dmmu0.page_table\[3\]\[1\] _0900_ vssd1 vssd1 vccd1
+ vccd1 _0951_ sky130_fd_sc_hd__mux2_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _2932_ dmmu1.page_table\[10\]\[6\] _2922_ _2933_ vssd1 vssd1 vccd1 vccd1 _0398_
+ sky130_fd_sc_hd__a31o_1
XFILLER_285_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5624__A1 _2240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7389__A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5029_ _2301_ immu_0.page_table\[15\]\[7\] _2298_ _2309_ vssd1 vssd1 vccd1 vccd1
+ _0782_ sky130_fd_sc_hd__a31o_1
XANTENNA__4806__A _2084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7059__CLK clknet_leaf_80_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5927__A2 _2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3938__A1 _1447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3856__S net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4541__A _1967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input273_A dcache_wb_sel[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6468__A _2190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5372__A _1944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4115__A1 _1584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5803__C _2750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4666__A2 _2083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5091__B _2338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3323__C1 _0906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6407__A3 _3116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3766__S _0839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4451__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6576__CLK clknet_leaf_46_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4400_ net325 net379 icache_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__mux2_1
XFILLER_145_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5380_ _1929_ _2440_ vssd1 vssd1 vccd1 vccd1 _2524_ sky130_fd_sc_hd__or2_1
XANTENNA__5551__B1 _2625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput505 net505 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[27] sky130_fd_sc_hd__buf_2
Xoutput516 net516 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[8] sky130_fd_sc_hd__buf_2
Xoutput527 net527 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[15] sky130_fd_sc_hd__buf_2
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4331_ _1831_ _1832_ _1833_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__nand3_1
Xoutput538 net538 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[3] sky130_fd_sc_hd__buf_2
Xoutput549 net549 vssd1 vssd1 vccd1 vccd1 dcache_mem_i_data[12] sky130_fd_sc_hd__buf_2
XFILLER_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7050_ clknet_leaf_36_core_clock _0311_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4262_ immu_1.page_table\[12\]\[8\] immu_1.page_table\[13\]\[8\] _1524_ vssd1 vssd1
+ vccd1 vccd1 _1768_ sky130_fd_sc_hd__mux2_1
XANTENNA__5713__C _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6001_ _2795_ _2881_ vssd1 vssd1 vccd1 vccd1 _2886_ sky130_fd_sc_hd__and2_1
X_3213_ _0827_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_1
X_4193_ immu_1.page_table\[12\]\[7\] immu_1.page_table\[13\]\[7\] _1443_ vssd1 vssd1
+ vccd1 vccd1 _1700_ sky130_fd_sc_hd__mux2_1
XANTENNA__3865__A0 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_23_core_clock_A clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_227_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3960__S0 _1472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6903_ clknet_leaf_76_core_clock _0164_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6834_ clknet_leaf_68_core_clock _0095_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6031__A1 _2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6919__CLK clknet_leaf_75_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6765_ clknet_leaf_85_core_clock _0026_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3977_ immu_1.page_table\[2\]\[1\] immu_1.page_table\[3\]\[1\] _1443_ vssd1 vssd1
+ vccd1 vccd1 _1490_ sky130_fd_sc_hd__mux2_1
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4999__C _2282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5457__A _2312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5716_ _2249_ _2699_ _2714_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__a21o_1
X_6696_ clknet_leaf_41_core_clock _0766_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5647_ _2227_ _2669_ _2674_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__a21o_1
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5578_ _2633_ vssd1 vssd1 vccd1 vccd1 _2634_ sky130_fd_sc_hd__buf_2
XFILLER_163_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6288__A _2784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4529_ net197 vssd1 vssd1 vccd1 vccd1 _1995_ sky130_fd_sc_hd__buf_6
XFILLER_49_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5192__A _2216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7248_ clknet_leaf_20_core_clock _0509_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5623__C _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout710 net211 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_16
XFILLER_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3856__A0 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7179_ clknet_leaf_33_core_clock _0440_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[8\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5920__A _2834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input119_A c1_o_mem_addr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6599__CLK clknet_leaf_56_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3586__S _1169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5367__A _2300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input390_A inner_wb_i_dat[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4271__A _1447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5086__B _2338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input84_A c0_sr_bus_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4210__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5830__A _2777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 c0_o_instr_long_addr[4] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_2
XFILLER_36_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4446__A _1933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6261__A1 _3042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4165__B _1663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_89_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4811__A2 _2172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3900_ immu_0.page_table\[4\]\[0\] immu_0.page_table\[5\]\[0\] immu_0.page_table\[6\]\[0\]
+ immu_0.page_table\[7\]\[0\] _1407_ net313 vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__mux4_1
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4880_ net78 _2213_ net77 net91 vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__or4b_2
XANTENNA__6013__A1 _2884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3831_ _1368_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3496__S _0881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5277__A _2458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6550_ clknet_leaf_51_core_clock _0620_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3762_ net136 net31 _1322_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__mux2_2
XFILLER_257_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4612__C _2049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5501_ net99 _2593_ vssd1 vssd1 vccd1 vccd1 _2597_ sky130_fd_sc_hd__and2_1
X_3693_ net121 _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__or2_1
X_6481_ _1569_ net255 _3171_ _1911_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__o211a_1
XANTENNA__7492__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5432_ _2546_ immu_0.page_table\[6\]\[10\] _2540_ _2554_ vssd1 vssd1 vccd1 vccd1
+ _0131_ sky130_fd_sc_hd__a31o_1
XFILLER_145_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5363_ _1935_ _2512_ vssd1 vssd1 vccd1 vccd1 _2515_ sky130_fd_sc_hd__and2_1
XFILLER_126_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7102_ clknet_leaf_30_core_clock _0363_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[13\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_259_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4314_ immu_1.page_table\[4\]\[9\] immu_1.page_table\[5\]\[9\] _1439_ vssd1 vssd1
+ vccd1 vccd1 _1819_ sky130_fd_sc_hd__mux2_1
XFILLER_273_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5294_ _2473_ dmmu0.page_table\[14\]\[9\] _2464_ vssd1 vssd1 vccd1 vccd1 _2475_ sky130_fd_sc_hd__and3_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5827__A1 _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4245_ immu_0.page_table\[14\]\[8\] immu_0.page_table\[15\]\[8\] _1480_ vssd1 vssd1
+ vccd1 vccd1 _1751_ sky130_fd_sc_hd__mux2_1
X_7033_ clknet_leaf_13_core_clock _0294_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4176_ net113 immu_1.high_addr_off\[3\] vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__nand2_1
XFILLER_82_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3260__A _0853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6741__CLK clknet_leaf_66_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4263__B1 _1516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6004__A1 _2884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6817_ clknet_leaf_59_core_clock _0078_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6290__B _3060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4803__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5187__A _2400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4110__S0 _1437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6891__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6748_ clknet_leaf_67_core_clock _0009_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[13\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6679_ clknet_leaf_56_core_clock _0749_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7247__CLK clknet_leaf_26_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_91_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_136_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4869__A2 _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5818__A1 _2232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5650__A _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6491__A1 _1977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input236_A dcache_wb_adr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4266__A _1584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6243__A1 _3026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input403_A inner_wb_i_dat[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5809__B dmmu0.page_table\[3\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5349__A3 _2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5097__A _1922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4205__S _1472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4021__A3 _1515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4309__A1 _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3517__C1 _0957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5544__B _2621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output455_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6614__CLK clknet_leaf_54_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4030_ _1424_ _1538_ _1540_ _1432_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__o211a_1
XFILLER_84_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3296__A1 _0881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4176__A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3391__S1 _0864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5981_ _2867_ dmmu1.page_table\[13\]\[9\] _2859_ _2872_ vssd1 vssd1 vccd1 vccd1 _0362_
+ sky130_fd_sc_hd__a31o_1
X_4932_ _2237_ dmmu0.page_table\[0\]\[12\] _2220_ vssd1 vssd1 vccd1 vccd1 _2254_ sky130_fd_sc_hd__and3_1
XANTENNA__4904__A _2204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6391__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4863_ _2182_ immu_1.page_table\[3\]\[5\] _2197_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__and3_1
XFILLER_220_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6602_ clknet_leaf_54_core_clock _0672_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[6\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3814_ _1358_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_1
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4794_ _2150_ immu_1.page_table\[4\]\[7\] _2157_ vssd1 vssd1 vccd1 vccd1 _2165_ sky130_fd_sc_hd__and3_1
X_6533_ clknet_leaf_45_core_clock _0603_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3745_ _0839_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__buf_4
XFILLER_158_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6464_ _2971_ immu_1.page_table\[8\]\[3\] _3159_ vssd1 vssd1 vccd1 vccd1 _3163_ sky130_fd_sc_hd__and3_1
X_3676_ _1255_ _1256_ _1257_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__and3_1
XFILLER_173_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5415_ _2531_ immu_0.page_table\[6\]\[2\] _2541_ _2545_ vssd1 vssd1 vccd1 vccd1 _0123_
+ sky130_fd_sc_hd__a31o_1
XFILLER_173_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6395_ net204 _3118_ vssd1 vssd1 vccd1 vccd1 _3123_ sky130_fd_sc_hd__and2_1
XANTENNA__5512__A3 _2591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5346_ _1944_ _2497_ vssd1 vssd1 vccd1 vccd1 _2505_ sky130_fd_sc_hd__and2_1
XFILLER_102_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5277_ _2458_ dmmu0.page_table\[14\]\[1\] _2464_ vssd1 vssd1 vccd1 vccd1 _2466_ sky130_fd_sc_hd__and3_1
XANTENNA__5470__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6473__A1 _1983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5276__A2 _2462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7016_ clknet_leaf_17_core_clock _0277_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[4\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4228_ _1732_ _1733_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__nor2_1
XANTENNA__6285__B _2153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4086__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4159_ _1584_ _1666_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__or2_1
XANTENNA__3382__S1 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7397__A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4787__A1 _2010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4814__A _2166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinterconnect_inner_720 vssd1 vssd1 vccd1 vccd1 interconnect_inner_720/HI c0_i_core_int_sreg[11]
+ sky130_fd_sc_hd__conb_1
XFILLER_184_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinterconnect_inner_731 vssd1 vssd1 vccd1 vccd1 interconnect_inner_731/HI c1_i_core_int_sreg[8]
+ sky130_fd_sc_hd__conb_1
XFILLER_7_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6637__CLK clknet_leaf_57_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input186_A c1_sr_bus_addr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input353_A ic1_mem_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6787__CLK clknet_leaf_0_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input47_A c0_o_mem_high_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6476__A _2190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5380__A _1929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6195__B _3002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3373__S1 _0864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4724__A _2121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4443__B _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5258__C _2445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput12 c0_o_instr_long_addr[7] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_2
XANTENNA__3774__S _0839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput23 c0_o_mem_addr[4] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 c0_o_mem_data[14] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
Xinput45 c0_o_mem_high_addr[0] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dlymetal6s2s_1
X_3530_ _1113_ _1114_ _0854_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__mux2_1
Xinput56 c0_o_mem_sel[1] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
Xinput67 c0_o_req_addr[2] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__buf_2
XFILLER_155_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput78 c0_sr_bus_addr[11] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_143_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput89 c0_sr_bus_addr[7] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
X_3461_ dmmu0.page_table\[14\]\[5\] dmmu0.page_table\[15\]\[5\] _0910_ vssd1 vssd1
+ vccd1 vccd1 _1049_ sky130_fd_sc_hd__mux2_1
XFILLER_170_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4163__C1 _1451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5200_ _2400_ dmmu0.page_table\[8\]\[3\] _2411_ vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__and3_1
XANTENNA__4702__A1 _2010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6180_ _2977_ dmmu1.page_table\[8\]\[9\] _2981_ _2993_ vssd1 vssd1 vccd1 vccd1 _0440_
+ sky130_fd_sc_hd__a31o_1
X_3392_ dmmu1.page_table\[4\]\[3\] dmmu1.page_table\[5\]\[3\] dmmu1.page_table\[6\]\[3\]
+ dmmu1.page_table\[7\]\[3\] _0858_ _0861_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__mux4_1
XFILLER_269_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5131_ _2211_ _2369_ _2374_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__a21o_1
XANTENNA__6386__A _3117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3803__A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5062_ _2316_ immu_0.page_table\[14\]\[8\] _2320_ _2330_ vssd1 vssd1 vccd1 vccd1
+ _0794_ sky130_fd_sc_hd__a31o_1
XFILLER_284_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4013_ immu_1.page_table\[14\]\[2\] immu_1.page_table\[15\]\[2\] _1524_ vssd1 vssd1
+ vccd1 vccd1 _1525_ sky130_fd_sc_hd__mux2_1
XFILLER_225_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4634__A _1999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4769__A1 _2021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5964_ _2805_ dmmu1.page_table\[13\]\[1\] _2859_ _2863_ vssd1 vssd1 vccd1 vccd1 _0354_
+ sky130_fd_sc_hd__a31o_1
XFILLER_252_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7092__CLK clknet_leaf_35_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5449__B _2559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4915_ net102 vssd1 vssd1 vccd1 vccd1 _2242_ sky130_fd_sc_hd__buf_6
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5895_ _2819_ dmmu0.page_table\[6\]\[7\] _2814_ vssd1 vssd1 vccd1 vccd1 _2823_ sky130_fd_sc_hd__and3_1
XANTENNA__5981__A3 _2859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5168__C _2392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4846_ _1987_ _2189_ _2192_ immu_1.page_table\[1\]\[9\] vssd1 vssd1 vccd1 vccd1 _0716_
+ sky130_fd_sc_hd__o22a_1
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3684__S _1146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4777_ _2154_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__clkbuf_4
XFILLER_165_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6516_ clknet_leaf_36_core_clock _0586_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3728_ _0854_ _1308_ net123 vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__a21oi_1
X_7496_ net398 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6447_ net213 net212 _0817_ _3152_ _1911_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__o311a_1
XFILLER_161_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3659_ _0901_ _1240_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__or2_1
XFILLER_134_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4154__C1 _1451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6378_ _3101_ dmmu1.page_table\[2\]\[11\] _3095_ _3111_ vssd1 vssd1 vccd1 vccd1 _0520_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5329_ _2494_ vssd1 vssd1 vccd1 vccd1 _2495_ sky130_fd_sc_hd__clkbuf_4
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6446__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5249__A2 _2442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3859__S net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4544__A _1972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6462__C _3159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input101_A c0_sr_bus_data_o[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5359__B _2512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3432__A1 _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_core_clock clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_98_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4719__A _2000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3623__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_28_core_clock_A clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4463__A3 _1924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4454__A _1898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4700_ _2008_ _2101_ _2108_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__a21o_1
XFILLER_187_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _2229_ immu_0.high_addr_off\[3\] _2690_ vssd1 vssd1 vccd1 vccd1 _2694_ sky130_fd_sc_hd__mux2_1
XFILLER_187_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4631_ _2062_ _2063_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__or2_2
XFILLER_187_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_68_core_clock clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__6952__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5285__A _2458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7350_ net304 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_2
X_4562_ _2019_ _2002_ _2020_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__a21o_1
XFILLER_265_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6301_ _3053_ dmmu1.page_table\[4\]\[5\] _3058_ _3066_ vssd1 vssd1 vccd1 vccd1 _0488_
+ sky130_fd_sc_hd__a31o_1
X_3513_ dmmu0.page_table\[12\]\[7\] dmmu0.page_table\[13\]\[7\] dmmu0.page_table\[14\]\[7\]
+ dmmu0.page_table\[15\]\[7\] _0896_ _0912_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__mux4_1
X_7281_ clknet_leaf_21_core_clock _0542_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4493_ _1967_ _1970_ vssd1 vssd1 vccd1 vccd1 _1971_ sky130_fd_sc_hd__and2_1
XFILLER_116_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7308__CLK clknet_leaf_19_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6232_ _3010_ dmmu1.page_table\[6\]\[3\] _3019_ _3025_ vssd1 vssd1 vccd1 vccd1 _0460_
+ sky130_fd_sc_hd__a31o_1
XFILLER_103_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3444_ _0881_ _1027_ _1031_ _0874_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__a211o_1
XFILLER_277_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6163_ _2791_ _2983_ vssd1 vssd1 vccd1 vccd1 _2985_ sky130_fd_sc_hd__and2_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3375_ _0964_ _0965_ _0887_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__mux2_1
XANTENNA__4629__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6428__A1 _3128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _1944_ _2355_ vssd1 vssd1 vccd1 vccd1 _2362_ sky130_fd_sc_hd__and2_1
XFILLER_257_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6094_ _1968_ _2099_ vssd1 vssd1 vccd1 vccd1 _2943_ sky130_fd_sc_hd__nor2_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5100__A1 _2347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5045_ _2316_ immu_0.page_table\[14\]\[0\] _2320_ _2321_ vssd1 vssd1 vccd1 vccd1
+ _0786_ sky130_fd_sc_hd__a31o_1
XFILLER_214_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5651__A2 _2669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4364__A _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6996_ clknet_leaf_6_core_clock _0257_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_240_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5947_ _2852_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5878_ _2443_ _2539_ vssd1 vssd1 vccd1 vccd1 _2813_ sky130_fd_sc_hd__or2_1
XANTENNA__5167__A1 _2227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5907__B _2555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4829_ _2182_ immu_1.page_table\[2\]\[10\] _2173_ vssd1 vssd1 vccd1 vccd1 _2186_
+ sky130_fd_sc_hd__and3_1
XFILLER_193_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_30_core_clock_A clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_166_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4914__A1 _2240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7479_ net176 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_2
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4539__A _1910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput202 c1_sr_bus_data_o[2] vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_2
Xinput213 dcache_mem_exception vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_2
XFILLER_102_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput224 dcache_mem_o_data[4] vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5890__A2 _2812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input149_A c1_o_mem_data[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput235 dcache_wb_adr[13] vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_2
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput246 dcache_wb_adr[23] vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_2
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput257 dcache_wb_o_dat[10] vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput268 dcache_wb_o_dat[6] vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_6
XFILLER_124_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput279 ic0_mem_data[11] vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_1
XFILLER_263_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6825__CLK clknet_leaf_59_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input316_A ic0_wb_adr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4274__A _1462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4705__C _2103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6198__A3 _3000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6975__CLK clknet_leaf_0_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4213__S _1407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4905__A1 _2233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6370__A3 _3096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput709 net709 vssd1 vssd1 vccd1 vccd1 inner_wb_we sky130_fd_sc_hd__buf_2
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4133__A2 _1636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4449__A _1935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5881__A2 _2812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3499__S _0872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4841__B1 _2192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6850_ clknet_leaf_70_core_clock _0111_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4615__C _2049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5801_ _2762_ dmmu0.page_table\[13\]\[11\] _2750_ vssd1 vssd1 vccd1 vccd1 _2764_
+ sky130_fd_sc_hd__and3_1
XANTENNA__5397__A1 _2531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6781_ clknet_leaf_86_core_clock _0042_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3993_ immu_0.page_table\[8\]\[2\] immu_0.page_table\[9\]\[2\] _1472_ vssd1 vssd1
+ vccd1 vccd1 _1505_ sky130_fd_sc_hd__mux2_2
XFILLER_62_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7495__A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5732_ immu_1.high_addr_off\[3\] _1974_ _2720_ vssd1 vssd1 vccd1 vccd1 _2724_ sky130_fd_sc_hd__mux2_1
XFILLER_222_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4912__A _2239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5149__A1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5663_ _2247_ _2669_ _2683_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__a21o_1
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7130__CLK clknet_leaf_29_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7402_ net341 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_1
XFILLER_148_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4614_ _1897_ vssd1 vssd1 vccd1 vccd1 _2054_ sky130_fd_sc_hd__buf_2
X_5594_ _2640_ dmmu0.page_table\[12\]\[7\] _2634_ vssd1 vssd1 vccd1 vccd1 _2643_ sky130_fd_sc_hd__and3_1
XANTENNA__4350__C _1411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4545_ _1910_ immu_1.page_table\[14\]\[2\] _2004_ vssd1 vssd1 vccd1 vccd1 _2009_
+ sky130_fd_sc_hd__and3_1
XFILLER_190_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5743__A _2729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7264_ clknet_leaf_19_core_clock _0525_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4476_ net194 net193 net192 net210 vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__or4b_1
XFILLER_89_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5462__B _2572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6215_ _3010_ dmmu1.page_table\[7\]\[10\] _2999_ _3014_ vssd1 vssd1 vccd1 vccd1 _0454_
+ sky130_fd_sc_hd__a31o_1
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5321__A1 _2489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3427_ dmmu0.page_table\[4\]\[4\] dmmu0.page_table\[5\]\[4\] dmmu0.page_table\[6\]\[4\]
+ dmmu0.page_table\[7\]\[4\] _0897_ _0902_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__mux4_1
X_7195_ clknet_leaf_27_core_clock _0456_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[7\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3263__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6848__CLK clknet_leaf_69_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5181__C _2392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _2971_ dmmu0.page_table\[1\]\[9\] _2962_ vssd1 vssd1 vccd1 vccd1 _2973_ sky130_fd_sc_hd__and3_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ dmmu0.page_table\[0\]\[1\] dmmu0.page_table\[1\]\[1\] _0910_ vssd1 vssd1 vccd1
+ vccd1 _0950_ sky130_fd_sc_hd__mux2_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _2801_ _2924_ vssd1 vssd1 vccd1 vccd1 _2933_ sky130_fd_sc_hd__and2_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3289_ dmmu1.page_table\[0\]\[0\] dmmu1.page_table\[1\]\[0\] _0865_ vssd1 vssd1 vccd1
+ vccd1 _0882_ sky130_fd_sc_hd__mux2_1
XFILLER_180_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5624__A2 _2650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5028_ _1944_ _2302_ vssd1 vssd1 vccd1 vccd1 _2309_ sky130_fd_sc_hd__and2_1
XANTENNA__6998__CLK clknet_leaf_39_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4806__B _2170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5388__A1 _2517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6979_ clknet_leaf_57_core_clock _0240_ vssd1 vssd1 vccd1 vccd1 immu_0.high_addr_off\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_241_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5918__A _2834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4822__A _2105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3494__S0 _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4348__C1 _1416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4033__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3872__S _1390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input266_A dcache_wb_o_dat[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6104__A3 _2942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5372__B _2512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4115__A2 _1623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5312__A1 _2363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7003__CLK clknet_leaf_36_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5379__A1 _2517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5828__A _2777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7153__CLK clknet_leaf_30_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4732__A _2121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output485_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5551__A1 _2229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput506 net506 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[28] sky130_fd_sc_hd__buf_2
Xoutput517 net517 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[9] sky130_fd_sc_hd__buf_2
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput528 net528 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[16] sky130_fd_sc_hd__buf_2
X_4330_ _1831_ _1832_ _1833_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__a21o_1
XFILLER_125_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput539 net539 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[4] sky130_fd_sc_hd__buf_2
XFILLER_125_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6500__A0 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4261_ _1523_ _1766_ vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__nor2_1
XFILLER_262_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6000_ _2884_ dmmu1.page_table\[12\]\[2\] _2878_ _2885_ vssd1 vssd1 vccd1 vccd1 _0368_
+ sky130_fd_sc_hd__a31o_1
X_3212_ net226 _0824_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__and2_1
XFILLER_79_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4192_ _1454_ _1696_ _1698_ _1451_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__o211a_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4907__A _2235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3960__S1 _1419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3811__A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6902_ clknet_leaf_79_core_clock _0163_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6833_ clknet_leaf_66_core_clock _0094_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_250_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4642__A _1897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6764_ clknet_leaf_87_core_clock _0025_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3976_ _1451_ _1488_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__or2_1
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6520__CLK clknet_leaf_43_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5457__B _2559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5715_ _2709_ dmmu0.page_table\[2\]\[10\] _2701_ vssd1 vssd1 vccd1 vccd1 _2714_ sky130_fd_sc_hd__and3_1
X_6695_ clknet_leaf_42_core_clock _0765_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3258__A _0852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5646_ _2666_ dmmu0.page_table\[11\]\[2\] _2671_ vssd1 vssd1 vccd1 vccd1 _2674_ sky130_fd_sc_hd__and3_1
XFILLER_108_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6334__A3 _3077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5542__A1 _2618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3692__S net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5577_ _2443_ _2334_ vssd1 vssd1 vccd1 vccd1 _2633_ sky130_fd_sc_hd__or2_1
XANTENNA__6670__CLK clknet_leaf_2_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4528_ _1976_ dmmu1.page_table\[14\]\[12\] _1963_ _1994_ vssd1 vssd1 vccd1 vccd1
+ _0596_ sky130_fd_sc_hd__a31o_1
XANTENNA__6288__B _2153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5192__B _2407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7247_ clknet_leaf_26_core_clock _0508_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[3\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4459_ _1942_ _1931_ vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__and2_1
XFILLER_277_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7026__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7178_ clknet_leaf_33_core_clock _0439_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[8\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_277_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3400__S0 _0898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3856__A1 _1381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ _2845_ dmmu0.page_table\[1\]\[1\] _2962_ vssd1 vssd1 vccd1 vccd1 _2964_ sky130_fd_sc_hd__and3_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7176__CLK clknet_leaf_34_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4028__S _1407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5648__A _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6470__C _3159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5230__B1 _2434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5781__A1 _2223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input383_A ic1_wb_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6325__A3 _3077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5533__A1 _2603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input77_A c0_sr_bus_addr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3631__A _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4446__B _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5064__A3 _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4272__A1 _1581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6543__CLK clknet_leaf_50_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3830_ _1363_ net266 vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__and2_1
XANTENNA__4462__A _1944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3761_ _1330_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_2
XANTENNA__5772__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6693__CLK clknet_leaf_43_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5500_ _2588_ immu_0.page_table\[3\]\[3\] _2591_ _2596_ vssd1 vssd1 vccd1 vccd1 _0157_
+ sky130_fd_sc_hd__a31o_1
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6480_ inner_wb_arbiter.o_sel_sig net255 _1899_ vssd1 vssd1 vccd1 vccd1 _3171_ sky130_fd_sc_hd__a21bo_1
XFILLER_158_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3692_ dmmu1.page_table\[4\]\[11\] dmmu1.page_table\[5\]\[11\] net120 vssd1 vssd1
+ vccd1 vccd1 _1274_ sky130_fd_sc_hd__mux2_1
XFILLER_200_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6316__A3 _3057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5431_ _2314_ _2543_ vssd1 vssd1 vccd1 vccd1 _2554_ sky130_fd_sc_hd__and2_1
XANTENNA__6389__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4401__S _0811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7049__CLK clknet_leaf_32_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5362_ _2503_ immu_0.page_table\[8\]\[2\] _2510_ _2514_ vssd1 vssd1 vccd1 vccd1 _0101_
+ sky130_fd_sc_hd__a31o_1
XFILLER_99_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7101_ clknet_leaf_31_core_clock _0362_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[13\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4313_ _1523_ _1815_ _1817_ _1530_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__o211a_1
XFILLER_141_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5293_ _2245_ _2462_ _2474_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__a21o_1
XFILLER_113_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7032_ clknet_leaf_13_core_clock _0293_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4244_ _1420_ _1749_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__or2_1
XFILLER_87_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4175_ _1596_ _1674_ _1677_ _1615_ vssd1 vssd1 vccd1 vccd1 _1682_ sky130_fd_sc_hd__o211a_1
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4263__A1 _1581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3687__S _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5468__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6816_ clknet_leaf_60_core_clock _0077_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5187__B dmmu0.page_table\[9\]\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4110__S1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6747_ clknet_leaf_66_core_clock _0008_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[13\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3959_ net312 vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__buf_6
XFILLER_167_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3774__A0 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6678_ clknet_leaf_55_core_clock _0748_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5629_ _2655_ dmmu0.page_table\[15\]\[9\] _2652_ vssd1 vssd1 vccd1 vccd1 _2663_ sky130_fd_sc_hd__and3_1
XANTENNA__5515__A1 _2603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4311__S _1438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4547__A _1974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input131_A c1_o_mem_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6566__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input229_A dcache_mem_o_data[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3597__S _1169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5378__A _2314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4713__C _2103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5097__B _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5754__A1 _2229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5506__A1 _2588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3612__S0 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output448_A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6909__CLK clknet_leaf_76_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5980_ _1987_ _2861_ vssd1 vssd1 vccd1 vccd1 _2872_ sky130_fd_sc_hd__and2_1
XFILLER_264_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4931_ net95 vssd1 vssd1 vccd1 vccd1 _2253_ sky130_fd_sc_hd__buf_4
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6391__B _3118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4862_ _1977_ _2195_ _2202_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__a21o_1
XFILLER_268_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4623__C _2049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6601_ clknet_leaf_54_core_clock _0671_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[6\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3813_ net220 _1348_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__and2_1
XFILLER_220_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4793_ _2016_ _2155_ _2164_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__a21o_1
XFILLER_220_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3756__A0 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6532_ clknet_leaf_46_core_clock _0602_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3744_ _1321_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4920__A _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6463_ _1972_ _3157_ _3162_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__a21o_1
XFILLER_173_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_35_core_clock_A clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_118_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3675_ net156 dmmu1.long_off_reg\[6\] vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__nand2_1
X_5414_ net97 _2543_ vssd1 vssd1 vccd1 vccd1 _2545_ sky130_fd_sc_hd__and2_1
XANTENNA__6170__A1 _2977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6394_ _3112_ dmmu1.page_table\[1\]\[3\] _3116_ _3122_ vssd1 vssd1 vccd1 vccd1 _0525_
+ sky130_fd_sc_hd__a31o_1
X_5345_ _2503_ immu_0.page_table\[9\]\[6\] _2495_ _2504_ vssd1 vssd1 vccd1 vccd1 _0094_
+ sky130_fd_sc_hd__a31o_1
XFILLER_141_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6589__CLK clknet_leaf_44_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5276_ _2211_ _2462_ _2465_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__a21o_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5470__B _2577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7015_ clknet_leaf_11_core_clock _0276_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[4\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6473__A2 _3157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4227_ net9 immu_0.high_addr_off\[4\] vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__nor2_1
XANTENNA__4367__A _1584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3271__A _0863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4158_ immu_1.page_table\[6\]\[6\] immu_1.page_table\[7\]\[6\] _1453_ vssd1 vssd1
+ vccd1 vccd1 _1666_ sky130_fd_sc_hd__mux2_1
XFILLER_233_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4086__B immu_1.high_addr_off\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4089_ _1569_ _1598_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__nor2_1
XFILLER_243_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4787__A2 _2155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3444__C1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5198__A _2400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4306__S _1524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5629__C _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5736__A1 _1979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinterconnect_inner_721 vssd1 vssd1 vccd1 vccd1 interconnect_inner_721/HI c0_i_core_int_sreg[12]
+ sky130_fd_sc_hd__conb_1
Xinterconnect_inner_732 vssd1 vssd1 vccd1 vccd1 interconnect_inner_732/HI c1_i_core_int_sreg[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5926__A _2834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_core_clock clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_194_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input179_A c1_o_req_addr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5661__A _2681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input346_A ic1_mem_data[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5380__B _2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4277__A net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5019__A3 _2298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5975__A1 _2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3986__A0 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_58_core_clock clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_187_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5836__A _1958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4740__A _2121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 c0_o_mem_addr[0] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput24 c0_o_mem_addr[5] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
Xinput35 c0_o_mem_data[15] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_155_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput46 c0_o_mem_high_addr[1] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
Xinput57 c0_o_mem_we vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3356__A _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput68 c0_o_req_addr[3] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_2
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput79 c0_sr_bus_addr[12] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
X_3460_ _0909_ _1045_ _1047_ _0918_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__o211a_1
XFILLER_182_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4702__A2 _2101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3391_ dmmu1.page_table\[0\]\[3\] dmmu1.page_table\[1\]\[3\] dmmu1.page_table\[2\]\[3\]
+ dmmu1.page_table\[3\]\[3\] _0892_ _0864_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__mux4_1
XFILLER_170_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5130_ _2371_ dmmu0.page_table\[10\]\[0\] _2373_ vssd1 vssd1 vccd1 vccd1 _2374_ sky130_fd_sc_hd__and3_1
XFILLER_69_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3803__B _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5061_ _2310_ _2322_ vssd1 vssd1 vccd1 vccd1 _2330_ sky130_fd_sc_hd__and2_1
XANTENNA__4187__A _1447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6881__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4466__A1 _1939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4012_ _1448_ vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__buf_6
XFILLER_272_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7498__A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4915__A net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5963_ _2791_ _2861_ vssd1 vssd1 vccd1 vccd1 _2863_ sky130_fd_sc_hd__and2_1
XANTENNA__4769__A2 _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5966__A1 _2805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4634__B _2064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5430__A3 _2541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4914_ _2240_ _2219_ _2241_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__a21o_1
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5894_ _2239_ _2812_ _2822_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__a21o_1
XFILLER_178_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4845_ _1985_ _2189_ _2192_ immu_1.page_table\[1\]\[8\] vssd1 vssd1 vccd1 vccd1 _0715_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__5718__A1 _2251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5746__A _2709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4776_ _2000_ _2153_ vssd1 vssd1 vccd1 vccd1 _2154_ sky130_fd_sc_hd__nor2_1
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6515_ clknet_leaf_43_core_clock _0585_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3727_ dmmu1.page_table\[4\]\[12\] dmmu1.page_table\[5\]\[12\] dmmu1.page_table\[6\]\[12\]
+ dmmu1.page_table\[7\]\[12\] _1146_ net121 vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__mux4_1
XFILLER_193_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7495_ net397 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3266__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6446_ net562 _3151_ mem_dcache_arb.select vssd1 vssd1 vccd1 vccd1 _3152_ sky130_fd_sc_hd__a21o_1
X_3658_ dmmu0.page_table\[8\]\[11\] dmmu0.page_table\[9\]\[11\] _0895_ vssd1 vssd1
+ vccd1 vccd1 _1240_ sky130_fd_sc_hd__mux2_1
XANTENNA__4629__B_N net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6377_ net199 _3097_ vssd1 vssd1 vccd1 vccd1 _3111_ sky130_fd_sc_hd__and2_1
X_3589_ _0901_ _1172_ _0905_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__a21oi_1
XFILLER_88_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5328_ _1929_ _2388_ vssd1 vssd1 vccd1 vccd1 _2494_ sky130_fd_sc_hd__or2_1
XFILLER_102_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6296__B _3060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5259_ _2243_ _2442_ _2454_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__a21o_1
XFILLER_244_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4457__A1 _1939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4825__A _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4036__S _1472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6604__CLK clknet_leaf_53_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3432__A2 _1006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3875__S _1390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5656__A _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4560__A _1983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input296_A ic0_mem_data[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6134__A1 _2229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4145__B1 _1360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5391__A _2300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4719__B _2118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_5_0_core_clock_A clknet_2_2_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5948__A1 _1937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4620__A1 _2016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4630_ net188 net181 vssd1 vssd1 vccd1 vccd1 _2063_ sky130_fd_sc_hd__nand2_1
XANTENNA__4470__A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4561_ _2017_ immu_1.page_table\[14\]\[7\] _2004_ vssd1 vssd1 vccd1 vccd1 _2020_
+ sky130_fd_sc_hd__and3_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6300_ net205 _3060_ vssd1 vssd1 vccd1 vccd1 _3066_ sky130_fd_sc_hd__and2_1
XFILLER_190_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3512_ _1096_ _1097_ _0918_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__mux2_1
XFILLER_265_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7280_ clknet_leaf_21_core_clock _0541_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4492_ _1969_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__buf_2
XFILLER_6_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6231_ _2795_ _3021_ vssd1 vssd1 vccd1 vccd1 _3025_ sky130_fd_sc_hd__and2_1
X_3443_ _0869_ _1028_ _1030_ _0855_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__o211a_1
XANTENNA__5479__A3 _2574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4687__A1 _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6162_ _2977_ dmmu1.page_table\[8\]\[0\] _2981_ _2984_ vssd1 vssd1 vccd1 vccd1 _0431_
+ sky130_fd_sc_hd__a31o_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ dmmu1.page_table\[8\]\[2\] dmmu1.page_table\[9\]\[2\] dmmu1.page_table\[10\]\[2\]
+ dmmu1.page_table\[11\]\[2\] _0892_ _0861_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__mux4_1
XFILLER_281_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _2347_ immu_0.page_table\[13\]\[6\] _2353_ _2361_ vssd1 vssd1 vccd1 vccd1
+ _0005_ sky130_fd_sc_hd__a31o_1
XFILLER_257_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6093_ _2941_ vssd1 vssd1 vccd1 vccd1 _2942_ sky130_fd_sc_hd__clkbuf_4
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _1926_ _2319_ vssd1 vssd1 vccd1 vccd1 _2321_ sky130_fd_sc_hd__nor2_1
XFILLER_257_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4645__A _2072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6627__CLK clknet_leaf_41_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6995_ clknet_leaf_1_core_clock _0256_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_253_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5403__A3 _2525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5179__C _2392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5946_ dmmu0.long_off_reg\[3\] _1935_ _2848_ vssd1 vssd1 vccd1 vccd1 _2852_ sky130_fd_sc_hd__mux2_1
XFILLER_230_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4611__A1 _2008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6777__CLK clknet_leaf_81_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5877_ _2811_ vssd1 vssd1 vccd1 vccd1 _2812_ sky130_fd_sc_hd__buf_4
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5476__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4828_ _2023_ _2172_ _2185_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__a21o_1
XANTENNA__6364__A1 _3101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5167__A2 _2390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4914__A2 _2219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4759_ _2010_ _2138_ _2144_ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__a21o_1
XFILLER_239_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6116__A1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7478_ net175 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__buf_2
XFILLER_107_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6429_ net205 _3137_ vssd1 vssd1 vccd1 vccd1 _3143_ sky130_fd_sc_hd__and2_1
XFILLER_68_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5642__C _2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_255_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6100__A _2793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3350__A1 _0869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput203 c1_sr_bus_data_o[3] vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_2
Xinput214 dcache_mem_o_data[0] vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_4
XFILLER_130_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput225 dcache_mem_o_data[5] vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_4
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput236 dcache_wb_adr[14] vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
XFILLER_88_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput247 dcache_wb_adr[2] vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_4
XFILLER_276_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput258 dcache_wb_o_dat[11] vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput269 dcache_wb_o_dat[7] vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_6
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input211_A core_reset vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4274__B _1770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input309_A ic0_wb_adr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3956__A3 immu_0.page_table\[15\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_9_core_clock clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6355__A1 _3085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4905__A2 _2219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7082__CLK clknet_leaf_5_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4449__B _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output430_A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output528_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5094__A1 _2347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4465__A _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4841__A1 _1977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5800_ _1950_ _2747_ _2763_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__a21o_1
X_6780_ clknet_leaf_89_core_clock _0041_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3992_ immu_0.page_table\[10\]\[2\] immu_0.page_table\[11\]\[2\] _1480_ vssd1 vssd1
+ vccd1 vccd1 _1504_ sky130_fd_sc_hd__mux2_1
XANTENNA__4054__C1 _1457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5731_ _2723_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5296__A _2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3809__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6346__A1 _3085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5662_ _2682_ dmmu0.page_table\[11\]\[9\] _2671_ vssd1 vssd1 vccd1 vccd1 _2683_ sky130_fd_sc_hd__and3_1
XANTENNA__5149__A2 _2369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7401_ net340 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_1
X_4613_ _2010_ _2047_ _2053_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__a21o_1
XFILLER_175_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5593_ _2240_ _2632_ _2642_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__a21o_1
XFILLER_209_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4544_ _1972_ vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__buf_6
XFILLER_116_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7263_ clknet_leaf_20_core_clock _0524_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4475_ net195 _1953_ net196 vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__or3b_4
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6214_ _2895_ _3001_ vssd1 vssd1 vccd1 vccd1 _3014_ sky130_fd_sc_hd__and2_1
XFILLER_171_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3426_ dmmu0.page_table\[0\]\[4\] dmmu0.page_table\[1\]\[4\] dmmu0.page_table\[2\]\[4\]
+ dmmu0.page_table\[3\]\[4\] _0897_ _0902_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__mux4_1
X_7194_ clknet_leaf_27_core_clock _0455_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[7\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_277_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _1946_ _2960_ _2972_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__a21o_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3357_ dmmu0.page_table\[4\]\[1\] dmmu0.page_table\[5\]\[1\] dmmu0.page_table\[6\]\[1\]
+ dmmu0.page_table\[7\]\[1\] _0898_ _0948_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__mux4_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6076_ _2931_ vssd1 vssd1 vccd1 vccd1 _2932_ sky130_fd_sc_hd__buf_4
XFILLER_218_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3288_ _0872_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__buf_4
XFILLER_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5085__A1 _2332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5027_ _2301_ immu_0.page_table\[15\]\[6\] _2298_ _2308_ vssd1 vssd1 vccd1 vccd1
+ _0781_ sky130_fd_sc_hd__a31o_1
XANTENNA__4375__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6978_ clknet_leaf_77_core_clock _0239_ vssd1 vssd1 vccd1 vccd1 immu_0.high_addr_off\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_241_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5929_ _1946_ _2830_ _2842_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__a21o_1
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3494__S1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4314__S _1439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5934__A _2681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6468__C _3159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input161_A c1_o_mem_sel[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input259_A dcache_wb_o_dat[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3323__A1 _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6942__CLK clknet_leaf_85_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input22_A c0_o_mem_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5828__B dmmu0.page_table\[3\]\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6005__A _2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4339__B1 _1535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5000__A1 _1983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5844__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5551__A2 _2623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput507 net507 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[29] sky130_fd_sc_hd__buf_2
Xoutput518 net518 vssd1 vssd1 vccd1 vccd1 c1_i_req_data_valid sky130_fd_sc_hd__buf_2
Xoutput529 net529 vssd1 vssd1 vccd1 vccd1 dcache_mem_addr[17] sky130_fd_sc_hd__buf_2
XANTENNA__3364__A _0929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4260_ immu_1.page_table\[14\]\[8\] immu_1.page_table\[15\]\[8\] _1524_ vssd1 vssd1
+ vccd1 vccd1 _1766_ sky130_fd_sc_hd__mux2_1
XFILLER_140_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3211_ _0826_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_1
X_4191_ _1446_ _1697_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__or2_1
XFILLER_67_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5067__A1 _2332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3811__B _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6901_ clknet_leaf_72_core_clock _0162_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_235_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6832_ clknet_leaf_68_core_clock _0093_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4923__A _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6031__A3 _2902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6763_ clknet_leaf_86_core_clock _0024_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3975_ immu_1.page_table\[4\]\[1\] immu_1.page_table\[5\]\[1\] immu_1.page_table\[6\]\[1\]
+ immu_1.page_table\[7\]\[1\] _1437_ net367 vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__mux4_1
XANTENNA__3539__A net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5714_ _2247_ _2700_ _2713_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__a21o_1
X_6694_ clknet_leaf_41_core_clock _0764_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5645_ _2224_ _2669_ _2673_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__a21o_1
XFILLER_191_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6815__CLK clknet_leaf_0_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5576_ _2631_ vssd1 vssd1 vccd1 vccd1 _2632_ sky130_fd_sc_hd__clkbuf_4
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4527_ _1993_ _1969_ vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__and2_1
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3274__A _0864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7246_ clknet_leaf_26_core_clock _0507_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[3\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_236_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4458_ net101 vssd1 vssd1 vccd1 vccd1 _1942_ sky130_fd_sc_hd__buf_6
XANTENNA__4089__B _1598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3409_ _0872_ _0997_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__or2_1
X_7177_ clknet_leaf_33_core_clock _0438_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_4389_ net275 _1890_ _0811_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__mux2_4
XFILLER_98_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3400__S1 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6128_ _2210_ _2960_ _2963_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__a21o_1
XANTENNA__5920__C _2832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5058__A1 _2316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6059_ _2920_ vssd1 vssd1 vccd1 vccd1 _2921_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_42_core_clock_A clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5230__A1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5230__B2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5781__A2 _2748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5664__A _2682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input376_A ic1_wb_adr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5297__A1 _2249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6261__A3 _3038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4009__C1 _1457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7270__CLK clknet_leaf_25_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6013__A3 _2878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4462__B _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6838__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5277__C _2464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3760_ net135 net30 _1322_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__mux2_2
XANTENNA__5772__A2 _2729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3691_ dmmu1.page_table\[6\]\[11\] dmmu1.page_table\[7\]\[11\] _0856_ vssd1 vssd1
+ vccd1 vccd1 _1273_ sky130_fd_sc_hd__mux2_1
XFILLER_187_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5430_ _2546_ immu_0.page_table\[6\]\[9\] _2541_ _2553_ vssd1 vssd1 vccd1 vccd1 _0130_
+ sky130_fd_sc_hd__a31o_1
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6389__B _3118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5361_ _1933_ _2512_ vssd1 vssd1 vccd1 vccd1 _2514_ sky130_fd_sc_hd__and2_1
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5724__D _2272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4312_ _1581_ _1816_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__or2_1
X_7100_ clknet_leaf_32_core_clock _0361_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[13\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5292_ _2473_ dmmu0.page_table\[14\]\[8\] _2464_ vssd1 vssd1 vccd1 vccd1 _2474_ sky130_fd_sc_hd__and3_1
XFILLER_99_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5288__A1 _2240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7031_ clknet_leaf_6_core_clock _0292_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[13\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_259_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4243_ immu_0.page_table\[12\]\[8\] immu_0.page_table\[13\]\[8\] _1480_ vssd1 vssd1
+ vccd1 vccd1 _1749_ sky130_fd_sc_hd__mux2_1
XFILLER_99_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3822__A _1363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4174_ _1569_ net240 _1654_ _1681_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__a22o_4
XFILLER_95_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4129__S _1601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5460__A1 _2562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4653__A _2072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5468__B _2577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6004__A3 _2878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6815_ clknet_leaf_0_core_clock _0076_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[14\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5212__A1 _2245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6746_ clknet_leaf_67_core_clock _0007_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[13\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3958_ _1467_ _1468_ net315 _1470_ vssd1 vssd1 vccd1 vccd1 _1471_ sky130_fd_sc_hd__o211a_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4971__B1 _2277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3889_ _1404_ vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_1
X_6677_ clknet_leaf_56_core_clock _0747_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5484__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5628_ _2245_ _2650_ _2662_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__a21o_1
XFILLER_164_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_opt_1_0_core_clock_A clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5559_ _1929_ _2212_ vssd1 vssd1 vccd1 vccd1 _2626_ sky130_fd_sc_hd__or2_1
XFILLER_191_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7229_ clknet_leaf_22_core_clock _0490_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7143__CLK clknet_leaf_29_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3732__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5650__C _2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7293__CLK clknet_leaf_43_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input124_A c1_o_mem_addr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6243__A3 _3019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5563__A1_N _1926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3878__S _1390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4563__A _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5378__B _2512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_48_core_clock clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5754__A2 _2730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5394__A _1940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3517__A1 _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3612__S1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4738__A _2121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_87_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6660__CLK clknet_leaf_7_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4930_ _2251_ _2218_ _2252_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__a21o_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4904__C _2221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4861_ _2182_ immu_1.page_table\[3\]\[4\] _2197_ vssd1 vssd1 vccd1 vccd1 _2202_ sky130_fd_sc_hd__and3_1
XFILLER_60_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6600_ clknet_leaf_56_core_clock _0670_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3812_ _1357_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_1
XFILLER_60_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4792_ _2150_ immu_1.page_table\[4\]\[6\] _2157_ vssd1 vssd1 vccd1 vccd1 _2164_ sky130_fd_sc_hd__and3_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6531_ clknet_leaf_45_core_clock _0601_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3743_ net142 net37 _0847_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__mux2_2
XFILLER_146_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3817__A _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6462_ _2971_ immu_1.page_table\[8\]\[2\] _3159_ vssd1 vssd1 vccd1 vccd1 _3162_ sky130_fd_sc_hd__and3_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3674_ net156 dmmu1.long_off_reg\[6\] vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__or2_1
XFILLER_284_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5413_ _2531_ immu_0.page_table\[6\]\[1\] _2541_ _2544_ vssd1 vssd1 vccd1 vccd1 _0122_
+ sky130_fd_sc_hd__a31o_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6393_ net203 _3118_ vssd1 vssd1 vccd1 vccd1 _3122_ sky130_fd_sc_hd__and2_1
XFILLER_217_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5344_ _1942_ _2497_ vssd1 vssd1 vccd1 vccd1 _2504_ sky130_fd_sc_hd__and2_1
XFILLER_161_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5275_ _2458_ dmmu0.page_table\[14\]\[0\] _2464_ vssd1 vssd1 vccd1 vccd1 _2465_ sky130_fd_sc_hd__and3_1
XFILLER_99_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4226_ net9 immu_0.high_addr_off\[4\] vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__and2_1
X_7014_ clknet_leaf_38_core_clock _0275_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[4\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_275_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4157_ _1581_ _1664_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__or2_1
XFILLER_228_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4088_ _1462_ _1588_ _1594_ _1597_ _1579_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__o311a_1
XANTENNA__3698__S _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4383__A net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4814__C _2174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3995__A1 _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinterconnect_inner_711 vssd1 vssd1 vccd1 vccd1 interconnect_inner_711/HI c0_i_core_int_sreg[2]
+ sky130_fd_sc_hd__conb_1
Xinterconnect_inner_722 vssd1 vssd1 vccd1 vccd1 interconnect_inner_722/HI c0_i_core_int_sreg[13]
+ sky130_fd_sc_hd__conb_1
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinterconnect_inner_733 vssd1 vssd1 vccd1 vccd1 interconnect_inner_733/HI c1_i_core_int_sreg[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6729_ clknet_leaf_66_core_clock _0799_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6103__A _2795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6533__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4558__A _2017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput690 net690 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[0] sky130_fd_sc_hd__buf_2
XANTENNA__6476__C _3159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input241_A dcache_wb_adr[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input339_A ic1_mem_data[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5424__A1 _2546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5389__A _1935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4293__A _1424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3401__S _0906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4724__C _2123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7039__CLK clknet_leaf_13_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 c0_o_mem_addr[10] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_168_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4232__S _1408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 c0_o_mem_addr[6] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_167_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput36 c0_o_mem_data[1] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
Xinput47 c0_o_mem_high_addr[2] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_155_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput58 c0_o_req_active vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_2
XFILLER_6_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput69 c0_o_req_addr[4] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__buf_2
XANTENNA_output460_A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output558_A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4163__A1 _1581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3390_ _0893_ _0979_ _0887_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__o21a_2
XFILLER_170_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4468__A _1948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5060_ _2316_ immu_0.page_table\[14\]\[7\] _2320_ _2329_ vssd1 vssd1 vccd1 vccd1
+ _0793_ sky130_fd_sc_hd__a31o_1
XFILLER_257_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5663__A1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4011_ _1447_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__buf_4
XFILLER_77_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5415__A1 _2531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5962_ _2805_ dmmu1.page_table\[13\]\[0\] _2859_ _2862_ vssd1 vssd1 vccd1 vccd1 _0353_
+ sky130_fd_sc_hd__a31o_1
XFILLER_18_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4913_ _2237_ dmmu0.page_table\[0\]\[6\] _2221_ vssd1 vssd1 vccd1 vccd1 _2241_ sky130_fd_sc_hd__and3_1
XFILLER_178_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5893_ _2819_ dmmu0.page_table\[6\]\[6\] _2814_ vssd1 vssd1 vccd1 vccd1 _2822_ sky130_fd_sc_hd__and3_1
XANTENNA__4931__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4844_ _1983_ _2189_ _2192_ immu_1.page_table\[1\]\[7\] vssd1 vssd1 vccd1 vccd1 _0714_
+ sky130_fd_sc_hd__o22a_1
XFILLER_221_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4775_ net188 net181 _2117_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__or3_4
XFILLER_119_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6514_ clknet_leaf_36_core_clock _0584_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3726_ _0869_ _1304_ _1306_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__o21ai_1
X_7494_ net396 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_1
XANTENNA__6556__CLK clknet_leaf_50_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6445_ net213 net212 vssd1 vssd1 vccd1 vccd1 _3151_ sky130_fd_sc_hd__nor2_1
X_3657_ dmmu0.page_table\[10\]\[11\] dmmu0.page_table\[11\]\[11\] _0896_ vssd1 vssd1
+ vccd1 vccd1 _1239_ sky130_fd_sc_hd__mux2_1
XFILLER_106_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4154__A1 _1584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6376_ _3101_ dmmu1.page_table\[2\]\[10\] _3095_ _3110_ vssd1 vssd1 vccd1 vccd1 _0519_
+ sky130_fd_sc_hd__a31o_1
X_3588_ dmmu0.page_table\[10\]\[9\] dmmu0.page_table\[11\]\[9\] _1169_ vssd1 vssd1
+ vccd1 vccd1 _1172_ sky130_fd_sc_hd__mux2_1
XFILLER_88_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5327_ _2489_ immu_0.page_table\[10\]\[10\] _2479_ _2493_ vssd1 vssd1 vccd1 vccd1
+ _0087_ sky130_fd_sc_hd__a31o_1
XFILLER_244_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5258_ _2447_ dmmu0.page_table\[7\]\[7\] _2445_ vssd1 vssd1 vccd1 vccd1 _2454_ sky130_fd_sc_hd__and3_1
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4209_ immu_0.page_table\[0\]\[7\] immu_0.page_table\[1\]\[7\] _1425_ vssd1 vssd1
+ vccd1 vccd1 _1716_ sky130_fd_sc_hd__mux2_1
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5189_ net83 net76 _1913_ vssd1 vssd1 vccd1 vccd1 _2407_ sky130_fd_sc_hd__or3_4
XANTENNA__3665__B1 _0929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3417__B1 _1005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3432__A3 _1007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5937__A _2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input191_A c1_sr_bus_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input289_A ic0_mem_data[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6134__A2 _2960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3891__S _1386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4145__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input52_A c0_o_mem_high_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4288__A _1424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5645__A1 _2224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3920__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6070__A1 _2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4620__A2 _2047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5847__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6579__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output675_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5285__C _2464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4560_ _1983_ vssd1 vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__clkbuf_8
XFILLER_128_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3511_ dmmu0.page_table\[0\]\[7\] dmmu0.page_table\[1\]\[7\] dmmu0.page_table\[2\]\[7\]
+ dmmu0.page_table\[3\]\[7\] _0897_ _0902_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__mux4_1
X_4491_ _1968_ _1961_ vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__nor2_1
XFILLER_183_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3442_ _0863_ _1029_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__or2_1
XFILLER_6_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6230_ _3010_ dmmu1.page_table\[6\]\[2\] _3019_ _3024_ vssd1 vssd1 vccd1 vccd1 _0459_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__6397__B _3118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6161_ _2879_ _2983_ vssd1 vssd1 vccd1 vccd1 _2984_ sky130_fd_sc_hd__and2_1
X_3373_ dmmu1.page_table\[0\]\[2\] dmmu1.page_table\[1\]\[2\] dmmu1.page_table\[2\]\[2\]
+ dmmu1.page_table\[3\]\[2\] _0892_ _0864_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__mux4_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _1942_ _2355_ vssd1 vssd1 vccd1 vccd1 _2361_ sky130_fd_sc_hd__and2_1
X_6092_ _2940_ vssd1 vssd1 vccd1 vccd1 _2941_ sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6428__A3 _3135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _2319_ vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__clkbuf_4
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5100__A3 _2353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4926__A _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3830__A _1363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4137__S _1601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6994_ clknet_leaf_4_core_clock _0255_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_230_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_47_core_clock_A clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_225_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5945_ _2851_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4611__A2 _2047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5757__A _2736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5876_ _2216_ _2539_ vssd1 vssd1 vccd1 vccd1 _2811_ sky130_fd_sc_hd__nor2_1
XFILLER_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5476__B _2577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4827_ _2182_ immu_1.page_table\[2\]\[9\] _2174_ vssd1 vssd1 vccd1 vccd1 _2185_ sky130_fd_sc_hd__and3_1
XFILLER_193_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4758_ _2134_ immu_1.page_table\[5\]\[3\] _2140_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__and3_1
XFILLER_193_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3709_ _0908_ _1289_ _0905_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__o21ai_1
XFILLER_174_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7477_ net174 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__buf_2
X_4689_ _2000_ _2099_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__nor2_1
XANTENNA__5492__A _1925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6428_ _3128_ dmmu1.page_table\[0\]\[4\] _3135_ _3142_ vssd1 vssd1 vccd1 vccd1 _0539_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__5875__A1 _2805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6100__B _2944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6359_ net202 _3098_ vssd1 vssd1 vccd1 vccd1 _3102_ sky130_fd_sc_hd__and2_1
XFILLER_68_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4539__C _2004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput204 c1_sr_bus_data_o[4] vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
XFILLER_276_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3981__S0 _1493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput215 dcache_mem_o_data[10] vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_4
XFILLER_76_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput226 dcache_mem_o_data[6] vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_4
XFILLER_124_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput237 dcache_wb_adr[15] vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_2
XFILLER_48_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput248 dcache_wb_adr[3] vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_4
Xinput259 dcache_wb_o_dat[12] vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3638__B1 _1220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3740__A _1319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6052__A1 _2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input204_A c1_sr_bus_data_o[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4063__A0 immu_0.page_table\[8\]\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6721__CLK clknet_leaf_63_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3187__A inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6871__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3915__A _1424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7227__CLK clknet_leaf_22_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5618__A1 _2230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3650__A _0901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6291__A1 _3053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4465__B _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4841__A2 _2189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6043__A1 _2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4054__B1 _1462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5397__A3 _2525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3991_ _1478_ _1500_ _1502_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__a21o_1
XFILLER_250_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5577__A _2443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4481__A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5730_ immu_1.high_addr_off\[2\] _1972_ _2720_ vssd1 vssd1 vccd1 vccd1 _2723_ sky130_fd_sc_hd__mux2_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3809__B _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5661_ _2681_ vssd1 vssd1 vccd1 vccd1 _2682_ sky130_fd_sc_hd__clkbuf_4
X_7400_ net339 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_1
X_4612_ _2038_ immu_1.page_table\[12\]\[3\] _2049_ vssd1 vssd1 vccd1 vccd1 _2053_
+ sky130_fd_sc_hd__and3_1
XFILLER_175_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5554__B1 _2625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5592_ _2640_ dmmu0.page_table\[12\]\[6\] _2634_ vssd1 vssd1 vccd1 vccd1 _2642_ sky130_fd_sc_hd__and3_1
XFILLER_175_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4543_ _2006_ _2002_ _2007_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__a21o_1
XFILLER_190_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7262_ clknet_leaf_25_core_clock _0523_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6201__A _2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4474_ net187 net186 _1952_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__or3_1
XFILLER_104_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6213_ _3010_ dmmu1.page_table\[7\]\[9\] _3000_ _3013_ vssd1 vssd1 vccd1 vccd1 _0453_
+ sky130_fd_sc_hd__a31o_1
XFILLER_89_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3425_ _0918_ _1013_ _0899_ vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__o21a_1
X_7193_ clknet_leaf_29_core_clock _0454_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[7\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5321__A3 _2480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3356_ _0913_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__buf_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _2971_ dmmu0.page_table\[1\]\[8\] _2962_ vssd1 vssd1 vccd1 vccd1 _2972_ sky130_fd_sc_hd__and3_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6075_ _1897_ vssd1 vssd1 vccd1 vccd1 _2931_ sky130_fd_sc_hd__buf_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ net106 net158 _0879_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__o21a_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6282__A1 _3053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _1942_ _2302_ vssd1 vssd1 vccd1 vccd1 _2308_ sky130_fd_sc_hd__and2_1
XANTENNA__6744__CLK clknet_leaf_66_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ clknet_leaf_11_core_clock _0238_ vssd1 vssd1 vccd1 vccd1 immu_0.high_addr_off\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4045__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5388__A3 _2525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4596__A1 _2021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5918__C _2832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5928_ _2834_ dmmu0.page_table\[5\]\[8\] _2832_ vssd1 vssd1 vccd1 vccd1 _2842_ sky130_fd_sc_hd__and3_1
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5859_ net206 vssd1 vssd1 vccd1 vccd1 _2801_ sky130_fd_sc_hd__buf_2
XFILLER_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4348__A1 _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6111__A _2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3859__A0 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5312__A3 _2480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input154_A c1_o_mem_high_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4566__A _1987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6273__A1 _3042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input321_A ic0_wb_adr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input15_A c0_o_mem_addr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4587__A1 _2012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4131__S0 _1601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4732__C _2123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6005__B _2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4339__A1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5000__A2 _2280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6617__CLK clknet_leaf_62_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4240__S _1480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput508 net508 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[2] sky130_fd_sc_hd__buf_2
XFILLER_176_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput519 net519 vssd1 vssd1 vccd1 vccd1 c1_rst sky130_fd_sc_hd__buf_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output540_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output638_A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5860__A _2801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3210_ net225 _0824_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__and2_1
XFILLER_140_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4190_ immu_1.page_table\[10\]\[7\] immu_1.page_table\[11\]\[7\] net366 vssd1 vssd1
+ vccd1 vccd1 _1697_ sky130_fd_sc_hd__mux2_1
XANTENNA__3945__S0 _1437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3380__A _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4275__B1 inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6900_ clknet_leaf_75_core_clock _0161_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_242_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6016__A1 _2884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6831_ clknet_leaf_68_core_clock _0092_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6762_ clknet_leaf_87_core_clock _0023_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3974_ _1451_ _1484_ _1486_ net369 vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__o211a_1
XFILLER_210_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5713_ _2709_ dmmu0.page_table\[2\]\[9\] _2702_ vssd1 vssd1 vccd1 vccd1 _2713_ sky130_fd_sc_hd__and3_1
XFILLER_148_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6693_ clknet_leaf_43_core_clock _0763_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5644_ _2666_ dmmu0.page_table\[11\]\[1\] _2671_ vssd1 vssd1 vccd1 vccd1 _2673_ sky130_fd_sc_hd__and3_1
XFILLER_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5575_ _2217_ _2334_ vssd1 vssd1 vccd1 vccd1 _2631_ sky130_fd_sc_hd__nor2_2
X_4526_ net200 vssd1 vssd1 vccd1 vccd1 _1993_ sky130_fd_sc_hd__buf_2
X_7245_ clknet_leaf_26_core_clock _0506_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4457_ _1939_ immu_0.page_table\[11\]\[5\] _1924_ _1941_ vssd1 vssd1 vccd1 vccd1
+ _0578_ sky130_fd_sc_hd__a31o_1
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3408_ dmmu1.page_table\[12\]\[4\] dmmu1.page_table\[13\]\[4\] dmmu1.page_table\[14\]\[4\]
+ dmmu1.page_table\[15\]\[4\] _0891_ _0860_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__mux4_1
XFILLER_277_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7176_ clknet_leaf_34_core_clock _0437_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4388_ net329 net383 _1390_ vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__mux2_2
XANTENNA__3710__C1 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input7_A c0_o_instr_long_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6127_ _2845_ dmmu0.page_table\[1\]\[0\] _2962_ vssd1 vssd1 vccd1 vccd1 _2963_ sky130_fd_sc_hd__and3_1
X_3339_ dmmu1.page_table\[14\]\[1\] dmmu1.page_table\[15\]\[1\] _0865_ vssd1 vssd1
+ vccd1 vccd1 _0931_ sky130_fd_sc_hd__mux2_1
XFILLER_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3290__A _0864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _2919_ _2081_ vssd1 vssd1 vccd1 vccd1 _2920_ sky130_fd_sc_hd__or2_1
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5009_ _1922_ _2296_ vssd1 vssd1 vccd1 vccd1 _2297_ sky130_fd_sc_hd__or2_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_core_clock clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_214_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5648__C _2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7072__CLK clknet_leaf_79_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5230__A2 _2433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5533__A3 _2607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3465__A _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4741__A1 _2021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input271_A dcache_wb_o_dat[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input369_A ic1_wb_adr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4296__A _1419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_77_core_clock clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_209_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7400__A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3480__A1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4235__S _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3690_ _0868_ _1271_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__or2_1
XFILLER_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5360_ _2503_ immu_0.page_table\[8\]\[1\] _2510_ _2513_ vssd1 vssd1 vccd1 vccd1 _0100_
+ sky130_fd_sc_hd__a31o_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4311_ immu_1.page_table\[8\]\[9\] immu_1.page_table\[9\]\[9\] _1438_ vssd1 vssd1
+ vccd1 vccd1 _1816_ sky130_fd_sc_hd__mux2_1
XFILLER_273_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5291_ _2370_ vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__4387__A1_N _1885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5590__A _2640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5288__A2 _2462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6485__A1 _1967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7030_ clknet_leaf_7_core_clock _0291_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[13\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_4242_ _1478_ _1745_ _1747_ _1535_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__o211a_1
XFILLER_113_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3822__B net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4173_ _0813_ _1673_ _1680_ net664 vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__o31a_2
XFILLER_274_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3314__S _0906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6237__A1 _3026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7095__CLK clknet_leaf_37_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6814_ clknet_leaf_88_core_clock _0075_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[14\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5212__A2 _2409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6745_ clknet_leaf_66_core_clock _0006_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3957_ _1416_ _1469_ vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__or2_1
XFILLER_51_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5765__A _2736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4971__A1 _1974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6676_ clknet_leaf_55_core_clock _0746_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3888_ net232 _1403_ _1386_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__mux2_4
XFILLER_129_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5484__B _2577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5627_ _2655_ dmmu0.page_table\[15\]\[8\] _2652_ vssd1 vssd1 vccd1 vccd1 _2662_ sky130_fd_sc_hd__and3_1
XANTENNA__6932__CLK clknet_leaf_57_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3285__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4184__C1 _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5558_ _1950_ _2622_ _2624_ immu_0.page_table\[1\]\[10\] vssd1 vssd1 vccd1 vccd1
+ _0186_ sky130_fd_sc_hd__o22a_1
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4509_ _1981_ _1970_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__and2_1
XFILLER_183_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5489_ net85 net84 _1912_ vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__or3_4
XFILLER_78_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7228_ clknet_leaf_22_core_clock _0489_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7159_ clknet_leaf_12_core_clock _0420_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_263_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5005__A _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6228__A1 _3010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input117_A c1_o_instr_long_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6400__A1 _3112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5394__B _2527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input82_A c0_sr_bus_addr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5506__A3 _2591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4714__A1 _2023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3517__A2 _1098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3922__C1 _1411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6467__A1 _1977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3923__A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_257_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6219__A1 _3010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4754__A _2134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6805__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4860_ _1974_ _2195_ _2201_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__a21o_1
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3811_ net219 _1348_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__and2_1
XANTENNA__6955__CLK clknet_leaf_85_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4791_ _2014_ _2155_ _2163_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__a21o_1
XFILLER_177_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5585__A _2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6530_ clknet_leaf_42_core_clock _0600_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3742_ _1320_ vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4953__A1 _1981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4920__C _2221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6461_ _1967_ _3157_ _3161_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__a21o_1
XFILLER_118_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3673_ _1207_ _1208_ _1205_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__o21ai_1
XFILLER_146_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5412_ net96 _2543_ vssd1 vssd1 vccd1 vccd1 _2544_ sky130_fd_sc_hd__and2_1
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6392_ _3112_ dmmu1.page_table\[1\]\[2\] _3116_ _3121_ vssd1 vssd1 vccd1 vccd1 _0524_
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6170__A3 _2981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5343_ _2300_ vssd1 vssd1 vccd1 vccd1 _2503_ sky130_fd_sc_hd__clkbuf_4
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4929__A _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5274_ _2463_ vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__clkbuf_4
X_7013_ clknet_leaf_37_core_clock _0274_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4225_ _1569_ net241 _1731_ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__a21bo_4
XFILLER_268_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4156_ immu_1.page_table\[4\]\[6\] immu_1.page_table\[5\]\[6\] _1438_ vssd1 vssd1
+ vccd1 vccd1 _1664_ sky130_fd_sc_hd__mux2_1
XFILLER_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4087_ _1440_ _1595_ _1596_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__or3b_1
XFILLER_283_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3444__A1 _0881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5198__C _2411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5197__A1 _2224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4989_ _2284_ immu_1.page_table\[15\]\[2\] _2282_ vssd1 vssd1 vccd1 vccd1 _2286_
+ sky130_fd_sc_hd__and3_1
XFILLER_211_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinterconnect_inner_712 vssd1 vssd1 vccd1 vccd1 interconnect_inner_712/HI c0_i_core_int_sreg[3]
+ sky130_fd_sc_hd__conb_1
XANTENNA__5495__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinterconnect_inner_723 vssd1 vssd1 vccd1 vccd1 interconnect_inner_723/HI c0_i_core_int_sreg[14]
+ sky130_fd_sc_hd__conb_1
X_6728_ clknet_3_2_0_core_clock _0798_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xinterconnect_inner_734 vssd1 vssd1 vccd1 vccd1 interconnect_inner_734/HI c1_i_core_int_sreg[11]
+ sky130_fd_sc_hd__conb_1
XFILLER_137_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5926__C _2832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6659_ clknet_leaf_8_core_clock _0729_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6103__B _2944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7110__CLK clknet_leaf_35_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_54_core_clock_A clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_278_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4558__B immu_1.page_table\[14\]\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput680 net680 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[23] sky130_fd_sc_hd__buf_2
XANTENNA__7260__CLK clknet_leaf_25_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput691 net691 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[10] sky130_fd_sc_hd__buf_2
XFILLER_278_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input234_A dcache_wb_adr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4574__A _2000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input401_A inner_wb_i_dat[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5389__B _2527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4293__B _1797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5975__A3 _2859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5188__A1 _2253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3918__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4740__C _2123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput15 c0_o_mem_addr[11] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_4
Xinput26 c0_o_mem_addr[7] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput37 c0_o_mem_data[2] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput48 c0_o_mem_high_addr[3] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
Xinput59 c0_o_req_addr[0] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__buf_2
XFILLER_155_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5360__A1 _2503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output453_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4468__B _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5663__A2 _2669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4466__A3 _1924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4010_ net369 _1517_ _1521_ _1441_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__o211a_1
XFILLER_284_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5961_ _1995_ _2861_ vssd1 vssd1 vccd1 vccd1 _2862_ sky130_fd_sc_hd__and2_1
XFILLER_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5966__A3 _2859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4912_ _2239_ vssd1 vssd1 vccd1 vccd1 _2240_ sky130_fd_sc_hd__buf_4
XFILLER_279_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5892_ _2235_ _2812_ _2821_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__a21o_1
X_4843_ _1981_ _2189_ _2192_ immu_1.page_table\[1\]\[6\] vssd1 vssd1 vccd1 vccd1 _0713_
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3828__A _1363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5746__C _2732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4774_ _2025_ _2137_ _2152_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__a21o_1
XFILLER_119_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6513_ clknet_leaf_60_core_clock _0583_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[11\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3725_ _0859_ _1305_ _0871_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__o21a_1
X_7493_ net389 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_1
X_6444_ _1898_ dmmu1.page_table\[0\]\[12\] _3134_ _3150_ vssd1 vssd1 vccd1 vccd1 _0547_
+ sky130_fd_sc_hd__a31o_1
XFILLER_228_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3656_ net18 _1233_ _1237_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__or3_1
XFILLER_134_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7283__CLK clknet_leaf_25_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4154__A2 _1659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5351__A1 _2503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6375_ net198 _3097_ vssd1 vssd1 vccd1 vccd1 _3110_ sky130_fd_sc_hd__and2_1
XFILLER_164_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3587_ _0909_ _1170_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__nand2_1
XFILLER_114_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_core_clock clknet_2_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
X_5326_ _2314_ _2482_ vssd1 vssd1 vccd1 vccd1 _2493_ sky130_fd_sc_hd__and2_1
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5103__A1 _2347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5257_ _2240_ _2442_ _2453_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__a21o_1
XFILLER_275_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4457__A3 _1924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4208_ _1430_ _1712_ _1714_ _1432_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__o211a_1
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5188_ _2253_ _2389_ _2406_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__a21o_1
XFILLER_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3665__A1 _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4139_ _1479_ _1642_ _1644_ _1646_ _1413_ vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__a221o_1
XFILLER_228_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4825__C _2174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3968__A2 immu_0.page_table\[8\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5656__C _2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input184_A c1_sr_bus_addr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5342__A1 _2489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4569__A _1989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6650__CLK clknet_leaf_39_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input351_A ic1_mem_data[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input45_A c0_o_mem_high_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5645__A2 _2669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7006__CLK clknet_leaf_80_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7156__CLK clknet_leaf_29_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4243__S _1480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5863__A _2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3510_ dmmu0.page_table\[4\]\[7\] dmmu0.page_table\[5\]\[7\] dmmu0.page_table\[6\]\[7\]
+ dmmu0.page_table\[7\]\[7\] _0897_ _0902_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__mux4_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4490_ _1958_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__clkbuf_4
XFILLER_6_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3441_ dmmu1.page_table\[12\]\[5\] dmmu1.page_table\[13\]\[5\] _0857_ vssd1 vssd1
+ vccd1 vccd1 _1029_ sky130_fd_sc_hd__mux2_1
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3344__B1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6160_ _2982_ vssd1 vssd1 vccd1 vccd1 _2983_ sky130_fd_sc_hd__buf_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _0893_ _0962_ _0855_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__o21a_2
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5111_ _2347_ immu_0.page_table\[13\]\[5\] _2353_ _2360_ vssd1 vssd1 vccd1 vccd1
+ _0004_ sky130_fd_sc_hd__a31o_1
XFILLER_88_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _2919_ _2099_ vssd1 vssd1 vccd1 vccd1 _2940_ sky130_fd_sc_hd__or2_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5042_ _1922_ _2318_ vssd1 vssd1 vccd1 vccd1 _2319_ sky130_fd_sc_hd__or2_1
XFILLER_97_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4844__B1 _2192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3830__B net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4645__C _2068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6993_ clknet_leaf_5_core_clock _0254_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5944_ dmmu0.long_off_reg\[2\] _1933_ _2848_ vssd1 vssd1 vccd1 vccd1 _2851_ sky130_fd_sc_hd__mux2_1
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6523__CLK clknet_leaf_44_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5875_ _2805_ dmmu1.page_table\[15\]\[12\] _2786_ _2810_ vssd1 vssd1 vccd1 vccd1
+ _0318_ sky130_fd_sc_hd__a31o_1
X_4826_ _2021_ _2172_ _2184_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__a21o_1
XFILLER_193_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6364__A3 _3096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5572__A1 _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4757_ _2008_ _2138_ _2143_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__a21o_1
XFILLER_239_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3992__S _1480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5773__A _2216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6673__CLK clknet_leaf_58_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3708_ dmmu0.page_table\[14\]\[12\] dmmu0.page_table\[15\]\[12\] _0895_ vssd1 vssd1
+ vccd1 vccd1 _1289_ sky130_fd_sc_hd__mux2_1
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7476_ net173 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__buf_2
XANTENNA__6116__A3 _2942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4688_ _2027_ _2062_ vssd1 vssd1 vccd1 vccd1 _2099_ sky130_fd_sc_hd__or2_4
XFILLER_111_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6427_ net204 _3137_ vssd1 vssd1 vccd1 vccd1 _3142_ sky130_fd_sc_hd__and2_1
XFILLER_108_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3639_ net50 dmmu0.long_off_reg\[5\] vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__nand2_1
XFILLER_108_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6358_ _1910_ vssd1 vssd1 vccd1 vccd1 _3101_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__7029__CLK clknet_leaf_7_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5309_ _1933_ _2482_ vssd1 vssd1 vccd1 vccd1 _2484_ sky130_fd_sc_hd__and2_1
XFILLER_142_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6289_ _3059_ vssd1 vssd1 vccd1 vccd1 _3060_ sky130_fd_sc_hd__buf_2
XANTENNA__3981__S1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput205 c1_sr_bus_data_o[5] vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_2
Xinput216 dcache_mem_o_data[11] vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_4
XFILLER_276_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput227 dcache_mem_o_data[7] vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_4
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput238 dcache_wb_adr[16] vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_2
XFILLER_124_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput249 dcache_wb_adr[4] vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_4
XFILLER_271_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3638__B2 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7179__CLK clknet_leaf_33_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6109__A _2801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5013__A _1897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3497__S0 _0891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input399_A inner_wb_i_dat[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6355__A3 _3096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7403__A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3931__A _1442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5618__A2 _2650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6546__CLK clknet_leaf_50_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4762__A _2134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3990_ _1419_ _1501_ net315 vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__a21o_1
XANTENNA__4054__A1 _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5577__B _2334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4481__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6696__CLK clknet_leaf_41_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5660_ _1896_ vssd1 vssd1 vccd1 vccd1 _2681_ sky130_fd_sc_hd__clkbuf_4
XFILLER_200_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4611_ _2008_ _2047_ _2052_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__a21o_1
XANTENNA__5554__A1 _2239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5591_ _2236_ _2632_ _2641_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__a21o_1
XFILLER_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4542_ _1910_ immu_1.page_table\[14\]\[1\] _2004_ vssd1 vssd1 vccd1 vccd1 _2007_
+ sky130_fd_sc_hd__and3_1
XFILLER_128_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_1_0_core_clock_A clknet_2_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_7261_ clknet_leaf_20_core_clock _0522_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4473_ net185 net184 net183 net182 vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__or4_1
XANTENNA__6201__B _3002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6212_ _2893_ _3002_ vssd1 vssd1 vccd1 vccd1 _3013_ sky130_fd_sc_hd__and2_1
X_3424_ dmmu0.page_table\[12\]\[4\] dmmu0.page_table\[13\]\[4\] dmmu0.page_table\[14\]\[4\]
+ dmmu0.page_table\[15\]\[4\] _0897_ _0913_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__mux4_1
XANTENNA__4002__A _1432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7192_ clknet_leaf_27_core_clock _0453_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[7\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3412__S0 _0865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _2681_ vssd1 vssd1 vccd1 vccd1 _2971_ sky130_fd_sc_hd__buf_6
XFILLER_258_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4937__A _2084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _0945_ _0946_ _0918_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__mux2_2
XFILLER_225_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3841__A _1373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _2914_ dmmu1.page_table\[10\]\[5\] _2922_ _2930_ vssd1 vssd1 vccd1 vccd1 _0397_
+ sky130_fd_sc_hd__a31o_1
XFILLER_218_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3286_ net158 _0878_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__nand2_4
XFILLER_273_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4148__S _1437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5085__A3 _2336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5025_ _2301_ immu_0.page_table\[15\]\[5\] _2298_ _2307_ vssd1 vssd1 vccd1 vccd1
+ _0780_ sky130_fd_sc_hd__a31o_1
XFILLER_273_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4672__A _2089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_core_clock clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4045__A1 _1448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6976_ clknet_leaf_78_core_clock _0237_ vssd1 vssd1 vccd1 vccd1 immu_0.high_addr_off\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4596__A2 _2030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5793__A1 _2242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5927_ _2242_ _2830_ _2841_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__a21o_1
XFILLER_241_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3288__A _0872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5858_ _2618_ dmmu1.page_table\[15\]\[5\] _2787_ _2800_ vssd1 vssd1 vccd1 vccd1 _0311_
+ sky130_fd_sc_hd__a31o_1
XFILLER_110_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4348__A2 _1849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4809_ _1996_ _2172_ _2175_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__a21o_1
X_5789_ _2235_ _2748_ _2757_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__a21o_1
XFILLER_119_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7459_ net398 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6111__B _2944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3859__A1 _1383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3751__A _1325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6569__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input147_A c1_o_mem_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_67_core_clock clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input314_A ic0_wb_adr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4582__A _2017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4587__A2 _2030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4131__S1 _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3198__A _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3926__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6302__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput509 net509 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[30] sky130_fd_sc_hd__buf_2
XFILLER_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5860__B _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output533_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3945__S1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4275__A1 _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6830_ clknet_leaf_68_core_clock _0091_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3600__S _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4923__C _2221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6761_ clknet_leaf_93_core_clock _0022_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[10\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_3973_ _1447_ net368 _1485_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__or3_1
XFILLER_195_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5712_ _2245_ _2700_ _2712_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__a21o_1
X_6692_ clknet_leaf_42_core_clock _0762_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5643_ _2211_ _2669_ _2672_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__a21o_1
XANTENNA__5527__A1 _2603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3836__A _1363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6212__A _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5574_ _1950_ _2626_ _2630_ immu_0.page_table\[0\]\[10\] vssd1 vssd1 vccd1 vccd1
+ _0197_ sky130_fd_sc_hd__o22a_1
XFILLER_117_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3633__S0 _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4525_ _1976_ dmmu1.page_table\[14\]\[11\] _1963_ _1992_ vssd1 vssd1 vccd1 vccd1
+ _0595_ sky130_fd_sc_hd__a31o_1
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7244_ clknet_leaf_23_core_clock _0505_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_4456_ _1940_ _1931_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__and2_1
XFILLER_104_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3407_ _0994_ _0876_ _0877_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__nor3_1
XANTENNA__4667__A _2072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7175_ clknet_leaf_11_core_clock _0436_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4387_ _1885_ _1889_ _1569_ net246 vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3571__A _0869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_59_core_clock_A clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6126_ _2961_ vssd1 vssd1 vccd1 vccd1 _2962_ sky130_fd_sc_hd__clkbuf_4
X_3338_ _0890_ _0894_ _0930_ _0819_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__o22a_2
XFILLER_105_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5058__A3 _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6057_ _1958_ vssd1 vssd1 vccd1 vccd1 _2919_ sky130_fd_sc_hd__buf_2
XFILLER_285_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ dmmu1.page_table\[12\]\[0\] dmmu1.page_table\[13\]\[0\] dmmu1.page_table\[14\]\[0\]
+ dmmu1.page_table\[15\]\[0\] _0858_ _0861_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__mux4_1
XFILLER_252_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6861__CLK clknet_leaf_70_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5008_ _1912_ _2295_ vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__or2_4
XFILLER_73_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7217__CLK clknet_leaf_28_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5766__A1 _1948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6959_ clknet_leaf_87_core_clock _0220_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[15\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4341__S _1425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5664__C _2670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4741__A2 _2120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5961__A _1995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input264_A dcache_wb_o_dat[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3481__A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4009__B2 _1447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_61_core_clock_A clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_232_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3768__A0 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output483_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3656__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6032__A _2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3615__S0 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6734__CLK clknet_leaf_66_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4310_ immu_1.page_table\[10\]\[9\] immu_1.page_table\[11\]\[9\] _1524_ vssd1 vssd1
+ vccd1 vccd1 _1815_ sky130_fd_sc_hd__mux2_1
XFILLER_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5290_ _2243_ _2462_ _2472_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__a21o_1
XFILLER_126_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4241_ _1420_ _1746_ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__or2_1
Xclkbuf_3_7_0_core_clock clknet_2_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
X_4172_ _1440_ _1679_ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__nor2_1
XFILLER_267_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6207__A _2931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4653__C _2068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6813_ clknet_leaf_1_core_clock _0074_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[14\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_251_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4950__A _2262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6744_ clknet_leaf_66_core_clock _0005_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3956_ immu_0.page_table\[12\]\[1\] immu_0.page_table\[13\]\[1\] immu_0.page_table\[14\]\[1\]
+ immu_0.page_table\[15\]\[1\] net312 net313 vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__mux4_1
XFILLER_50_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6675_ clknet_leaf_56_core_clock _0745_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3887_ net310 net364 _1390_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__mux2_1
XANTENNA__4971__A2 _2274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3566__A _0868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4161__S _1437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5626_ _2243_ _2650_ _2661_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__a21o_1
XFILLER_176_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5557_ _1948_ _2623_ _2625_ immu_0.page_table\[1\]\[9\] vssd1 vssd1 vccd1 vccd1 _0185_
+ sky130_fd_sc_hd__o22a_1
XFILLER_247_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4508_ net206 vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__buf_6
XFILLER_132_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5488_ _2561_ vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__clkbuf_4
XFILLER_117_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7227_ clknet_leaf_22_core_clock _0488_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4397__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4439_ net96 vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__buf_6
XFILLER_263_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5684__A0 _2235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7158_ clknet_leaf_12_core_clock _0419_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3695__C1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6109_ _2801_ _2944_ vssd1 vssd1 vccd1 vccd1 _2952_ sky130_fd_sc_hd__and2_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7089_ clknet_leaf_2_core_clock _0350_ vssd1 vssd1 vccd1 vccd1 dmmu0.long_off_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_219_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7501__A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5987__A1 _2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4336__S _1480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6607__CLK clknet_leaf_53_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6117__A _2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3240__S _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__A _2784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input381_A ic1_wb_sel[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6164__A1 _2977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3195__B _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input75_A c0_o_req_ppl_submit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4714__A2 _2101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6467__A2 _3157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4738__C _2123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4100__A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3686__C1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7411__A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3438__C1 _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4650__A1 _2016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5866__A _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3810_ _1356_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4770__A _2105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4790_ _2150_ immu_1.page_table\[4\]\[5\] _2157_ vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__and3_1
XFILLER_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3741_ net141 net36 _0847_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__mux2_1
XANTENNA__4953__A2 _2257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6460_ _2971_ immu_1.page_table\[8\]\[1\] _3159_ vssd1 vssd1 vccd1 vccd1 _3161_ sky130_fd_sc_hd__and3_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3672_ _1238_ _1247_ _1253_ _0957_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__a22o_1
XFILLER_185_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5411_ _1930_ _2539_ vssd1 vssd1 vccd1 vccd1 _2543_ sky130_fd_sc_hd__nor2_4
XFILLER_118_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5902__A1 _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6391_ net202 _3118_ vssd1 vssd1 vccd1 vccd1 _3121_ sky130_fd_sc_hd__and2_1
XFILLER_133_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5342_ _2489_ immu_0.page_table\[9\]\[5\] _2495_ _2502_ vssd1 vssd1 vccd1 vccd1 _0093_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__3913__B1 _1416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5273_ _2443_ _2318_ vssd1 vssd1 vccd1 vccd1 _2463_ sky130_fd_sc_hd__or2_1
XFILLER_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4469__A1 _1939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5106__A _1935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7012_ clknet_leaf_78_core_clock _0273_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4224_ inner_wb_arbiter.o_sel_sig _1706_ _1730_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__or3b_1
XANTENNA__7062__CLK clknet_leaf_10_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4155_ _1457_ _1658_ _1662_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__or3_1
XFILLER_233_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4086_ net110 immu_1.high_addr_off\[0\] vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__nand2_1
XFILLER_270_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4156__S _1438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4641__A1 _2008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5776__A _2443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4680__A _2089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5197__A2 _2409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6394__A1 _3112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4988_ _1967_ _2280_ _2285_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__a21o_1
XFILLER_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5495__B _2593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinterconnect_inner_713 vssd1 vssd1 vccd1 vccd1 interconnect_inner_713/HI c0_i_core_int_sreg[4]
+ sky130_fd_sc_hd__conb_1
X_6727_ clknet_leaf_66_core_clock _0797_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xinterconnect_inner_724 vssd1 vssd1 vccd1 vccd1 interconnect_inner_724/HI c0_i_core_int_sreg[15]
+ sky130_fd_sc_hd__conb_1
Xinterconnect_inner_735 vssd1 vssd1 vccd1 vccd1 interconnect_inner_735/HI c1_i_core_int_sreg[12]
+ sky130_fd_sc_hd__conb_1
X_3939_ _1437_ vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__buf_6
XFILLER_109_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6658_ clknet_leaf_43_core_clock _0728_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5609_ _2651_ vssd1 vssd1 vccd1 vccd1 _2652_ sky130_fd_sc_hd__buf_2
XFILLER_194_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6589_ clknet_leaf_44_core_clock _0659_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput670 net670 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[14] sky130_fd_sc_hd__buf_2
XFILLER_120_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput681 net681 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[2] sky130_fd_sc_hd__buf_2
XANTENNA__4558__C _2004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5016__A _1928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput692 net692 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[11] sky130_fd_sc_hd__buf_2
XFILLER_78_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4855__A _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input227_A dcache_mem_o_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4574__B _2028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5424__A3 _2541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput16 c0_o_mem_addr[12] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_4
XFILLER_128_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput27 c0_o_mem_addr[8] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4148__A0 immu_1.page_table\[14\]\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput38 c0_o_mem_data[3] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
Xinput49 c0_o_mem_high_addr[4] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3934__A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7406__A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7085__CLK clknet_leaf_93_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5360__A2 immu_0.page_table\[8\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output446_A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4871__A1 _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5415__A3 _2541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5960_ _2860_ vssd1 vssd1 vccd1 vccd1 _2861_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__4084__C1 _1553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4911_ net101 vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__buf_6
XFILLER_52_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5891_ _2819_ dmmu0.page_table\[6\]\[5\] _2814_ vssd1 vssd1 vccd1 vccd1 _2821_ sky130_fd_sc_hd__and3_1
XANTENNA__5596__A _2640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6376__A1 _3101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4842_ _1979_ _2189_ _2192_ immu_1.page_table\[1\]\[5\] vssd1 vssd1 vccd1 vccd1 _0712_
+ sky130_fd_sc_hd__o22a_1
XFILLER_20_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3828__B net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4773_ _2150_ immu_1.page_table\[5\]\[10\] _2139_ vssd1 vssd1 vccd1 vccd1 _2152_
+ sky130_fd_sc_hd__and3_1
XFILLER_165_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3724_ dmmu1.page_table\[0\]\[12\] dmmu1.page_table\[1\]\[12\] _1146_ vssd1 vssd1
+ vccd1 vccd1 _1305_ sky130_fd_sc_hd__mux2_1
X_6512_ clknet_leaf_58_core_clock _0582_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[11\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6128__A1 _2210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7492_ net211 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_1
XFILLER_228_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6443_ net200 _3136_ vssd1 vssd1 vccd1 vccd1 _3150_ sky130_fd_sc_hd__and2_1
X_3655_ _0908_ _1234_ _1236_ _0905_ vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__o211a_1
XANTENNA__3844__A _1375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6220__A _2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6374_ _3101_ dmmu1.page_table\[2\]\[9\] _3096_ _3109_ vssd1 vssd1 vccd1 vccd1 _0518_
+ sky130_fd_sc_hd__a31o_1
X_3586_ dmmu0.page_table\[8\]\[9\] dmmu0.page_table\[9\]\[9\] _1169_ vssd1 vssd1 vccd1
+ vccd1 _1170_ sky130_fd_sc_hd__mux2_1
XANTENNA__3362__A1 _0906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5325_ _2489_ immu_0.page_table\[10\]\[9\] _2480_ _2492_ vssd1 vssd1 vccd1 vccd1
+ _0086_ sky130_fd_sc_hd__a31o_1
XFILLER_248_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5256_ _2447_ dmmu0.page_table\[7\]\[6\] _2445_ vssd1 vssd1 vccd1 vccd1 _2453_ sky130_fd_sc_hd__and3_1
XFILLER_275_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4207_ _1423_ _1713_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__or2_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5187_ _2400_ dmmu0.page_table\[9\]\[12\] _2391_ vssd1 vssd1 vccd1 vccd1 _2406_ sky130_fd_sc_hd__and3_1
XANTENNA__4862__A1 _1977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4138_ _1570_ _1645_ _1535_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__o21a_1
XFILLER_244_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4069_ _0812_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__buf_4
XFILLER_260_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3968__A3 immu_0.page_table\[9\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4090__A2 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input177_A c1_o_req_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5342__A2 immu_0.page_table\[9\]\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input344_A ic1_mem_data[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6945__CLK clknet_leaf_85_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input38_A c0_o_mem_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6070__A3 _2922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3929__A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4369__B1 _1553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5863__B _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3440_ dmmu1.page_table\[14\]\[5\] dmmu1.page_table\[15\]\[5\] _0865_ vssd1 vssd1
+ vccd1 vccd1 _1028_ sky130_fd_sc_hd__mux2_1
XANTENNA__6040__A _2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3344__A1 _0872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3371_ _0960_ _0961_ _0887_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__mux2_1
XFILLER_124_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _1940_ _2355_ vssd1 vssd1 vccd1 vccd1 _2360_ sky130_fd_sc_hd__and2_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _2932_ dmmu1.page_table\[10\]\[12\] _2921_ _2939_ vssd1 vssd1 vccd1 vccd1
+ _0404_ sky130_fd_sc_hd__a31o_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _2295_ _2317_ vssd1 vssd1 vccd1 vccd1 _2318_ sky130_fd_sc_hd__or2_4
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4495__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4844__A1 _1983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7100__CLK clknet_leaf_32_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6992_ clknet_leaf_9_core_clock _0253_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_18_core_clock clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_280_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5943_ _2850_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_280_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5757__C _2732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5874_ _1993_ _2788_ vssd1 vssd1 vccd1 vccd1 _2810_ sky130_fd_sc_hd__and2_1
XANTENNA__3280__B1 _0872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4825_ _2182_ immu_1.page_table\[2\]\[8\] _2174_ vssd1 vssd1 vccd1 vccd1 _2184_ sky130_fd_sc_hd__and3_1
XANTENNA__5021__A1 _2301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6818__CLK clknet_leaf_59_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4756_ _2134_ immu_1.page_table\[5\]\[2\] _2140_ vssd1 vssd1 vccd1 vccd1 _2143_ sky130_fd_sc_hd__and3_1
XFILLER_146_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5773__B _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3707_ _0901_ _1287_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__nor2_1
XFILLER_119_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4687_ _2025_ _2082_ _2098_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__a21o_1
X_7475_ net172 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_2
X_3638_ _1215_ _1217_ _1220_ net18 vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__o22a_1
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6426_ _3128_ dmmu1.page_table\[0\]\[3\] _3135_ _3141_ vssd1 vssd1 vccd1 vccd1 _0538_
+ sky130_fd_sc_hd__a31o_1
XFILLER_104_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0_1_core_clock clknet_1_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_1_0_1_core_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_161_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3569_ _1145_ _1148_ _1150_ _1152_ net123 vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__o221a_2
X_6357_ _3085_ dmmu1.page_table\[2\]\[1\] _3096_ _3100_ vssd1 vssd1 vccd1 vccd1 _0510_
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5308_ _2363_ immu_0.page_table\[10\]\[1\] _2480_ _2483_ vssd1 vssd1 vccd1 vccd1
+ _0078_ sky130_fd_sc_hd__a31o_1
XFILLER_276_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6288_ _2784_ _2153_ vssd1 vssd1 vccd1 vccd1 _3059_ sky130_fd_sc_hd__nor2_2
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput206 c1_sr_bus_data_o[6] vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
XFILLER_88_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_core_clock clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_core_clock
+ sky130_fd_sc_hd__clkbuf_16
Xinput217 dcache_mem_o_data[12] vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_4
XFILLER_276_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput228 dcache_mem_o_data[8] vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput239 dcache_wb_adr[17] vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_2
X_5239_ _2441_ vssd1 vssd1 vccd1 vccd1 _2442_ sky130_fd_sc_hd__clkbuf_4
XFILLER_124_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6109__B _2944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4048__C1 _1441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3497__S1 _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3749__A _1324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6125__A _2215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_66_core_clock_A clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5012__A1 _1976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input294_A ic0_mem_data[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4220__C1 _1416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5079__A1 _2332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7123__CLK clknet_leaf_13_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4826__A1 _2021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6291__A3 _3058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output409_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7273__CLK clknet_leaf_26_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6043__A3 _2902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5251__A1 _2230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4054__A2 _1564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3659__A _0901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output680_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5874__A _1993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4610_ _2038_ immu_1.page_table\[12\]\[2\] _2049_ vssd1 vssd1 vccd1 vccd1 _2052_
+ sky130_fd_sc_hd__and3_1
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5590_ _2640_ dmmu0.page_table\[12\]\[5\] _2634_ vssd1 vssd1 vccd1 vccd1 _2641_ sky130_fd_sc_hd__and3_1
XANTENNA__5554__A2 _2623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4541_ _1967_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__buf_4
XFILLER_144_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7260_ clknet_leaf_25_core_clock _0521_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_4472_ _1939_ immu_0.page_table\[11\]\[10\] _1923_ _1951_ vssd1 vssd1 vccd1 vccd1
+ _0583_ sky130_fd_sc_hd__a31o_1
XFILLER_171_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6211_ _3010_ dmmu1.page_table\[7\]\[8\] _3000_ _3012_ vssd1 vssd1 vccd1 vccd1 _0452_
+ sky130_fd_sc_hd__a31o_1
X_3423_ _0906_ _1011_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__or2_1
X_7191_ clknet_leaf_28_core_clock _0452_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[7\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4002__B _1410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3412__S1 _0863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _2242_ _2960_ _2970_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__a21o_1
X_3354_ dmmu0.page_table\[8\]\[1\] dmmu0.page_table\[9\]\[1\] dmmu0.page_table\[10\]\[1\]
+ dmmu0.page_table\[11\]\[1\] _0910_ _0913_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__mux4_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4937__B _2255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _2799_ _2924_ vssd1 vssd1 vccd1 vccd1 _2930_ sky130_fd_sc_hd__and2_1
XFILLER_285_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3285_ net124 _0876_ _0877_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__or3_2
XFILLER_225_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__A1 _2012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5114__A _1944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _1940_ _2302_ vssd1 vssd1 vccd1 vccd1 _2307_ sky130_fd_sc_hd__and2_1
XFILLER_273_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6975_ clknet_leaf_0_core_clock _0236_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[11\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3253__A0 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5926_ _2834_ dmmu0.page_table\[5\]\[7\] _2832_ vssd1 vssd1 vccd1 vccd1 _2841_ sky130_fd_sc_hd__and3_1
XANTENNA__6640__CLK clknet_leaf_57_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5793__A2 _2748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5857_ _2799_ _2789_ vssd1 vssd1 vccd1 vccd1 _2800_ sky130_fd_sc_hd__and2_1
XFILLER_139_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5784__A _2749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4808_ _2166_ immu_1.page_table\[2\]\[0\] _2174_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__and3_1
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5788_ _2749_ dmmu0.page_table\[13\]\[5\] _2751_ vssd1 vssd1 vccd1 vccd1 _2757_ sky130_fd_sc_hd__and3_1
XFILLER_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6790__CLK clknet_leaf_80_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4739_ _2019_ _2120_ _2131_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__a21o_1
XFILLER_135_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7458_ net397 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_1
XFILLER_119_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6409_ _3128_ dmmu1.page_table\[1\]\[10\] _3115_ _3130_ vssd1 vssd1 vccd1 vccd1 _0532_
+ sky130_fd_sc_hd__a31o_1
XFILLER_1_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7389_ net359 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_1
XFILLER_162_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7504__A net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5024__A _1940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7296__CLK clknet_leaf_44_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6273__A3 _3038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5481__A1 _2576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5959__A _1968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4863__A _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3492__B1 _1078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input307_A ic0_mem_data[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5233__A1 _2223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3479__A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3244__A0 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5694__A _2682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6302__B _3060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3942__A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7414__A net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output526_A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4773__A _2150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6663__CLK clknet_leaf_9_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6016__A3 _2878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6760_ clknet_leaf_0_core_clock _0021_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[10\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3972_ immu_1.page_table\[10\]\[1\] immu_1.page_table\[11\]\[1\] _1443_ vssd1 vssd1
+ vccd1 vccd1 _1485_ sky130_fd_sc_hd__mux2_1
XFILLER_250_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7019__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5711_ _2709_ dmmu0.page_table\[2\]\[8\] _2702_ vssd1 vssd1 vccd1 vccd1 _2712_ sky130_fd_sc_hd__and3_1
XFILLER_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6691_ clknet_leaf_39_core_clock _0761_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5642_ _2666_ dmmu0.page_table\[11\]\[0\] _2671_ vssd1 vssd1 vccd1 vccd1 _2672_ sky130_fd_sc_hd__and3_1
XFILLER_176_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3836__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6212__B _3002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5573_ _1948_ _2627_ _2630_ immu_0.page_table\[0\]\[9\] vssd1 vssd1 vccd1 vccd1 _0196_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3633__S1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4524_ _1991_ _1969_ vssd1 vssd1 vccd1 vccd1 _1992_ sky130_fd_sc_hd__and2_1
XFILLER_144_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7243_ clknet_leaf_23_core_clock _0504_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4455_ net100 vssd1 vssd1 vccd1 vccd1 _1940_ sky130_fd_sc_hd__buf_6
XANTENNA__4948__A _2262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3852__A _1379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3406_ net106 _0994_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__and2_1
X_7174_ clknet_leaf_35_core_clock _0435_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4386_ net2 _1887_ _1888_ inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 _1889_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__3710__A1 _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3337_ _0898_ _0923_ _0929_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__mux2_1
X_6125_ _2215_ _2621_ vssd1 vssd1 vccd1 vccd1 _2961_ sky130_fd_sc_hd__or2_1
XFILLER_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_core_clock clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_258_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6056_ _2914_ dmmu1.page_table\[11\]\[12\] _2901_ _2918_ vssd1 vssd1 vccd1 vccd1
+ _0391_ sky130_fd_sc_hd__a31o_1
XFILLER_218_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3268_ _0860_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__buf_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3998__S _1408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ net85 net84 vssd1 vssd1 vccd1 vccd1 _2295_ sky130_fd_sc_hd__nand2_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3199_ net214 _0819_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__and2_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3299__A _0891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6958_ clknet_leaf_85_core_clock _0219_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[15\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5766__A2 _2730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4974__B1 _2277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5909_ _2443_ _2555_ vssd1 vssd1 vccd1 vccd1 _2831_ sky130_fd_sc_hd__or2_1
X_6889_ clknet_leaf_83_core_clock _0150_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6403__A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3238__S _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6536__CLK clknet_leaf_44_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5961__B _2861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3388__S0 _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input257_A dcache_wb_o_dat[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6686__CLK clknet_leaf_56_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5454__A1 _2562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A c0_o_mem_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4593__A _2038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5206__A1 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7409__A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7311__CLK clknet_leaf_2_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6313__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6032__B _2904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3615__S1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4768__A _2134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5590__C _2634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4240_ immu_0.page_table\[8\]\[8\] immu_0.page_table\[9\]\[8\] _1480_ vssd1 vssd1
+ vccd1 vccd1 _1746_ sky130_fd_sc_hd__mux2_1
XANTENNA__3379__S0 _0898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4487__B _1963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4171_ _1675_ _1678_ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__xor2_1
XFILLER_206_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6237__A3 _3019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3551__S0 _0897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6812_ clknet_leaf_87_core_clock _0073_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[14\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6743_ clknet_leaf_67_core_clock _0004_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3955_ immu_0.page_table\[10\]\[1\] immu_0.page_table\[11\]\[1\] _1425_ vssd1 vssd1
+ vccd1 vccd1 _1468_ sky130_fd_sc_hd__mux2_1
XFILLER_211_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3847__A _1373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6223__A _1968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5765__C _2732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6674_ clknet_leaf_58_core_clock _0744_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3886_ _1402_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__clkbuf_1
XANTENNA__6559__CLK clknet_leaf_48_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5625_ _2655_ dmmu0.page_table\[15\]\[7\] _2652_ vssd1 vssd1 vccd1 vccd1 _2661_ sky130_fd_sc_hd__and3_1
XFILLER_176_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4184__A1 _1523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5556_ _1946_ _2623_ _2625_ immu_0.page_table\[1\]\[8\] vssd1 vssd1 vccd1 vccd1 _0184_
+ sky130_fd_sc_hd__o22a_1
XFILLER_129_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4507_ _1976_ dmmu1.page_table\[14\]\[5\] _1964_ _1980_ vssd1 vssd1 vccd1 vccd1 _0589_
+ sky130_fd_sc_hd__a31o_1
XFILLER_2_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4678__A _2089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5487_ _2576_ immu_0.page_table\[4\]\[10\] _2573_ _2587_ vssd1 vssd1 vccd1 vccd1
+ _0153_ sky130_fd_sc_hd__a31o_1
XFILLER_172_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7226_ clknet_leaf_22_core_clock _0487_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4438_ _1911_ immu_0.page_table\[11\]\[0\] _1924_ _1927_ vssd1 vssd1 vccd1 vccd1
+ _0573_ sky130_fd_sc_hd__a31o_1
XFILLER_116_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7157_ clknet_leaf_13_core_clock _0418_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4369_ _1516_ _1866_ _1868_ _1553_ _1872_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__a311o_1
XFILLER_219_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6228__A3 _3019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6108_ _2948_ dmmu1.page_table\[9\]\[5\] _2942_ _2951_ vssd1 vssd1 vccd1 vccd1 _0410_
+ sky130_fd_sc_hd__a31o_1
XFILLER_112_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7088_ clknet_leaf_2_core_clock _0349_ vssd1 vssd1 vccd1 vccd1 dmmu0.long_off_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_246_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6039_ _2898_ dmmu1.page_table\[11\]\[4\] _2902_ _2909_ vssd1 vssd1 vccd1 vccd1 _0383_
+ sky130_fd_sc_hd__a31o_1
XFILLER_273_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5302__A _1922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__B _2028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6400__A3 _3116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3757__A _1328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4352__S _1524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6133__A _2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5972__A _2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input374_A ic1_wb_adr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4588__A _1897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input68_A c0_o_req_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4754__C _2140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5866__B _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6701__CLK clknet_leaf_42_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4262__S _1524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3740_ _1319_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5585__C _2634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3671_ _1249_ _1252_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__xnor2_1
XFILLER_118_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5882__A _2777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5410_ _2531_ immu_0.page_table\[6\]\[0\] _2541_ _2542_ vssd1 vssd1 vccd1 vccd1 _0121_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__6851__CLK clknet_leaf_69_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6390_ _3112_ dmmu1.page_table\[1\]\[1\] _3116_ _3120_ vssd1 vssd1 vccd1 vccd1 _0523_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__3913__A1 _1424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5341_ _1940_ _2497_ vssd1 vssd1 vccd1 vccd1 _2502_ sky130_fd_sc_hd__and2_1
XFILLER_154_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5272_ _2461_ vssd1 vssd1 vccd1 vccd1 _2462_ sky130_fd_sc_hd__buf_4
XANTENNA__7207__CLK clknet_leaf_27_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5106__B _2355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7011_ clknet_leaf_78_core_clock _0272_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4223_ net2 _1710_ _1711_ _1729_ _0812_ vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__a311o_1
X_4154_ _1584_ _1659_ _1661_ _1451_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__o211a_1
XFILLER_255_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5418__A1 _2546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6218__A _1993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_255_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3429__B1 _1017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4085_ net110 immu_1.high_addr_off\[0\] vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__nor2_1
XFILLER_283_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5776__B _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4987_ _2284_ immu_1.page_table\[15\]\[1\] _2282_ vssd1 vssd1 vccd1 vccd1 _2285_
+ sky130_fd_sc_hd__and3_1
XFILLER_168_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinterconnect_inner_714 vssd1 vssd1 vccd1 vccd1 interconnect_inner_714/HI c0_i_core_int_sreg[5]
+ sky130_fd_sc_hd__conb_1
X_6726_ clknet_leaf_61_core_clock _0796_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[14\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3601__B1 _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3938_ _1447_ _1449_ _1451_ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__a21o_1
XFILLER_211_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinterconnect_inner_725 vssd1 vssd1 vccd1 vccd1 interconnect_inner_725/HI c1_i_core_int_sreg[2]
+ sky130_fd_sc_hd__conb_1
XFILLER_258_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinterconnect_inner_736 vssd1 vssd1 vccd1 vccd1 interconnect_inner_736/HI c1_i_core_int_sreg[13]
+ sky130_fd_sc_hd__conb_1
XFILLER_183_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6657_ clknet_leaf_42_core_clock _0727_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3869_ net319 net373 _1390_ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__mux2_2
XFILLER_258_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5792__A _2749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5608_ _2443_ _2296_ vssd1 vssd1 vccd1 vccd1 _2651_ sky130_fd_sc_hd__or2_1
XFILLER_137_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6588_ clknet_leaf_45_core_clock _0658_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5539_ net104 _2609_ vssd1 vssd1 vccd1 vccd1 _2619_ sky130_fd_sc_hd__and2_1
XFILLER_127_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4201__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput660 net660 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[7] sky130_fd_sc_hd__buf_2
XANTENNA__5657__A1 _2243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput671 net671 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[15] sky130_fd_sc_hd__buf_2
XFILLER_160_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput682 net682 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[3] sky130_fd_sc_hd__buf_2
XANTENNA__5016__B _2302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7209_ clknet_leaf_15_core_clock _0470_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput693 net693 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[12] sky130_fd_sc_hd__buf_2
XFILLER_266_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3251__S _0847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6082__A1 _2932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input122_A c1_o_mem_addr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5967__A _2795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6874__CLK clknet_leaf_70_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 c0_o_mem_addr[13] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_2
Xinput28 c0_o_mem_addr[9] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput39 c0_o_mem_data[4] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3778__A_N net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5896__A1 _2242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5360__A3 _2510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5207__A _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4111__A _1619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output439_A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7422__A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_73_core_clock_A clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_237_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4871__A2 _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6038__A _2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5820__A1 _2235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4910_ _2236_ _2219_ _2238_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__a21o_1
XFILLER_280_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5890_ _2232_ _2812_ _2820_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__a21o_1
XFILLER_233_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4841_ _1977_ _2189_ _2192_ immu_1.page_table\[1\]\[4\] vssd1 vssd1 vccd1 vccd1 _0711_
+ sky130_fd_sc_hd__o22a_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4387__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4772_ _2023_ _2138_ _2151_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__a21o_1
XFILLER_165_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6511_ clknet_leaf_59_core_clock _0581_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[11\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3723_ dmmu1.page_table\[2\]\[12\] dmmu1.page_table\[3\]\[12\] _0857_ vssd1 vssd1
+ vccd1 vccd1 _1304_ sky130_fd_sc_hd__mux2_1
XFILLER_20_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7491_ net163 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_1
XANTENNA__6128__A2 _2960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4139__A1 _1479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6442_ _1898_ dmmu1.page_table\[0\]\[11\] _3134_ _3149_ vssd1 vssd1 vccd1 vccd1 _0546_
+ sky130_fd_sc_hd__a31o_1
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3654_ _0901_ _1235_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__or2_1
XANTENNA__6501__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5887__A1 _2229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6220__B _2118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6373_ net209 _3098_ vssd1 vssd1 vccd1 vccd1 _3109_ sky130_fd_sc_hd__and2_1
XANTENNA__5351__A3 _2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3585_ net15 vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__buf_6
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5117__A _2310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5324_ _2312_ _2482_ vssd1 vssd1 vccd1 vccd1 _2492_ sky130_fd_sc_hd__and2_1
XFILLER_161_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_47_core_clock clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_102_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4956__A _2262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5255_ _2236_ _2442_ _2452_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__a21o_1
XFILLER_275_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5103__A3 _2353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3860__A _1384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4206_ immu_0.page_table\[6\]\[7\] immu_0.page_table\[7\]\[7\] net312 vssd1 vssd1
+ vccd1 vccd1 _1713_ sky130_fd_sc_hd__mux2_1
XFILLER_275_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5186_ _2251_ _2389_ _2405_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__a21o_1
XANTENNA__6747__CLK clknet_leaf_66_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4862__A2 _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ immu_0.page_table\[0\]\[6\] immu_0.page_table\[1\]\[6\] _1601_ vssd1 vssd1
+ vccd1 vccd1 _1645_ sky130_fd_sc_hd__mux2_1
XFILLER_83_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6064__A1 _2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4068_ _1576_ _1577_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__nor2_1
XFILLER_209_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4691__A _2084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6897__CLK clknet_leaf_75_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4378__A1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6709_ clknet_leaf_63_core_clock _0779_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5726__S _2720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7507__A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_86_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5342__A3 _2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3246__S _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4866__A _2204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput490 net490 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[13] sky130_fd_sc_hd__buf_2
XFILLER_266_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input337_A ic1_mem_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5802__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4369__A1 _1516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4106__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7052__CLK clknet_leaf_32_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7417__A clknet_leaf_92_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5869__A1 _2805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output556_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6040__B _2904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3370_ dmmu1.page_table\[12\]\[2\] dmmu1.page_table\[13\]\[2\] dmmu1.page_table\[14\]\[2\]
+ dmmu1.page_table\[15\]\[2\] _0892_ _0864_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__mux4_1
XANTENNA__3975__S0 _1437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4776__A _2000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3727__S0 _1146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5040_ net76 net83 vssd1 vssd1 vccd1 vccd1 _2317_ sky130_fd_sc_hd__or2b_1
XFILLER_69_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3501__C1 _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4844__A2 _2189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4057__A0 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6991_ clknet_leaf_9_core_clock _0252_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_230_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5942_ dmmu0.long_off_reg\[1\] _1928_ _2848_ vssd1 vssd1 vccd1 vccd1 _2850_ sky130_fd_sc_hd__mux2_1
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5400__A _2310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5873_ _2805_ dmmu1.page_table\[15\]\[11\] _2786_ _2809_ vssd1 vssd1 vccd1 vccd1
+ _0317_ sky130_fd_sc_hd__a31o_1
XFILLER_240_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3280__A1 _0869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4824_ _2019_ _2172_ _2183_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__a21o_1
XANTENNA__5557__B1 _2625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4755_ _2006_ _2138_ _2142_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__a21o_1
XFILLER_159_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3706_ dmmu0.page_table\[12\]\[12\] dmmu0.page_table\[13\]\[12\] _1169_ vssd1 vssd1
+ vccd1 vccd1 _1287_ sky130_fd_sc_hd__mux2_1
XANTENNA__6231__A _2795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7474_ net171 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_1
X_4686_ _2089_ immu_1.page_table\[10\]\[10\] _2085_ vssd1 vssd1 vccd1 vccd1 _2098_
+ sky130_fd_sc_hd__and3_1
XFILLER_107_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6425_ net203 _3137_ vssd1 vssd1 vccd1 vccd1 _3141_ sky130_fd_sc_hd__and2_1
X_3637_ _1218_ _1219_ net17 vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__mux2_1
XFILLER_174_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6356_ net201 _3098_ vssd1 vssd1 vccd1 vccd1 _3100_ sky130_fd_sc_hd__and2_1
X_3568_ _0859_ _1151_ _0854_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__a21o_1
XFILLER_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5307_ _1928_ _2482_ vssd1 vssd1 vccd1 vccd1 _2483_ sky130_fd_sc_hd__and2_1
XANTENNA__4686__A _2089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6287_ _3057_ vssd1 vssd1 vccd1 vccd1 _3058_ sky130_fd_sc_hd__clkbuf_4
XFILLER_142_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3499_ _1083_ _1084_ _0872_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__mux2_1
Xinput207 c1_sr_bus_data_o[7] vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput218 dcache_mem_o_data[13] vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_4
XFILLER_76_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput229 dcache_mem_o_data[9] vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_4
X_5238_ _2217_ _2440_ vssd1 vssd1 vccd1 vccd1 _2441_ sky130_fd_sc_hd__nor2_1
XFILLER_276_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5169_ _2230_ _2390_ _2396_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__a21o_1
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6037__A1 _2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6406__A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7075__CLK clknet_leaf_10_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6125__B _2621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5548__B1 _2625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3765__A _1332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_1_0_core_clock clknet_1_0_1_core_clock vssd1 vssd1 vccd1 vccd1 clknet_2_1_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__6141__A _2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input287_A ic0_mem_data[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5980__A _1987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input50_A c0_o_mem_high_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4826__A2 _2172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4134__S0 _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4762__C _2140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5251__A2 _2442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6200__A1 _2994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output673_A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3675__A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4270__S _1437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6051__A _2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4540_ _1996_ _2002_ _2005_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__a21o_1
XFILLER_156_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6592__CLK clknet_leaf_44_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4471_ _1950_ _1931_ vssd1 vssd1 vccd1 vccd1 _1951_ sky130_fd_sc_hd__and2_1
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6210_ _2891_ _3002_ vssd1 vssd1 vccd1 vccd1 _3012_ sky130_fd_sc_hd__and2_1
X_3422_ dmmu0.page_table\[8\]\[4\] dmmu0.page_table\[9\]\[4\] dmmu0.page_table\[10\]\[4\]
+ dmmu0.page_table\[11\]\[4\] _0897_ _0913_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__mux4_1
X_7190_ clknet_leaf_15_core_clock _0451_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _2845_ dmmu0.page_table\[1\]\[7\] _2962_ vssd1 vssd1 vccd1 vccd1 _2970_ sky130_fd_sc_hd__and3_1
X_3353_ dmmu0.page_table\[12\]\[1\] dmmu0.page_table\[13\]\[1\] dmmu0.page_table\[14\]\[1\]
+ dmmu0.page_table\[15\]\[1\] _0910_ _0913_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__mux4_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3614__S net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6267__A1 _3042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6072_ _2914_ dmmu1.page_table\[10\]\[4\] _2922_ _2929_ vssd1 vssd1 vccd1 vccd1 _0396_
+ sky130_fd_sc_hd__a31o_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ net151 net150 net153 net152 vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__or4_1
XFILLER_258_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__A2 _2172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5114__B _2355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5023_ _2301_ immu_0.page_table\[15\]\[4\] _2298_ _2306_ vssd1 vssd1 vccd1 vccd1
+ _0779_ sky130_fd_sc_hd__a31o_1
XFILLER_285_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6019__A1 _2884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7098__CLK clknet_leaf_35_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_281_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6974_ clknet_leaf_0_core_clock _0235_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[11\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4672__C _2086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5130__A _2371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5925_ _2239_ _2830_ _2840_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__a21o_1
XFILLER_241_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5856_ net205 vssd1 vssd1 vccd1 vccd1 _2799_ sky130_fd_sc_hd__buf_2
XFILLER_194_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4807_ _2173_ vssd1 vssd1 vccd1 vccd1 _2174_ sky130_fd_sc_hd__buf_2
XANTENNA__6935__CLK clknet_leaf_58_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5787_ _2232_ _2748_ _2756_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__a21o_1
XFILLER_194_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3585__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4753__A1 _1996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4738_ _2121_ immu_1.page_table\[6\]\[7\] _2123_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__and3_1
XFILLER_5_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7457_ net396 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__clkbuf_1
XFILLER_119_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4669_ _1897_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__buf_2
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6408_ net198 _3117_ vssd1 vssd1 vccd1 vccd1 _3130_ sky130_fd_sc_hd__and2_1
XFILLER_102_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7388_ net358 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6339_ _2891_ _3079_ vssd1 vssd1 vccd1 vccd1 _3089_ sky130_fd_sc_hd__and2_1
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6258__A1 _3026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5024__B _2302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5959__B _2028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3492__A1 _0929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3492__B2 _0957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4582__C _2032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6430__A1 _3128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input202_A c1_sr_bus_data_o[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4992__A1 _1974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input98_A c0_sr_bus_data_o[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6497__A1 _1983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_12_core_clock_A clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_69_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3434__S _0865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6249__A1 _3026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5215__A _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6808__CLK clknet_leaf_85_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7430__A net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4265__S _1453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6046__A _2891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6958__CLK clknet_leaf_85_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3971_ immu_1.page_table\[12\]\[1\] immu_1.page_table\[13\]\[1\] immu_1.page_table\[14\]\[1\]
+ immu_1.page_table\[15\]\[1\] _1453_ _1454_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__mux4_1
XFILLER_211_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5710_ _2243_ _2700_ _2711_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__a21o_1
XFILLER_250_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6690_ clknet_leaf_58_core_clock _0760_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5641_ _2670_ vssd1 vssd1 vccd1 vccd1 _2671_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5527__A3 _2607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4196__C1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4735__A1 _2014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5572_ _1946_ _2627_ _2630_ immu_0.page_table\[0\]\[8\] vssd1 vssd1 vccd1 vccd1 _0195_
+ sky130_fd_sc_hd__o22a_1
X_7311_ clknet_leaf_2_core_clock _0572_ vssd1 vssd1 vccd1 vccd1 icore_sregs.c1_disable
+ sky130_fd_sc_hd__dfxtp_1
X_4523_ net199 vssd1 vssd1 vccd1 vccd1 _1991_ sky130_fd_sc_hd__buf_2
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7242_ clknet_leaf_21_core_clock _0503_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_4454_ _1898_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__buf_4
XFILLER_132_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3405_ net158 vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__inv_2
X_7173_ clknet_leaf_12_core_clock _0434_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4385_ _1831_ _1835_ _1886_ _1360_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__a31oi_1
XANTENNA__4667__C _2086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6124_ _2959_ vssd1 vssd1 vccd1 vccd1 _2960_ sky130_fd_sc_hd__clkbuf_4
X_3336_ _0927_ _0928_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__nor2_4
XFILLER_252_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _1993_ _2903_ vssd1 vssd1 vccd1 vccd1 _2918_ sky130_fd_sc_hd__and2_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _0859_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__buf_4
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _1989_ _2279_ _2294_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__a21o_1
XFILLER_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3198_ _0818_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__clkbuf_4
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ clknet_leaf_81_core_clock _0218_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4974__A1 _1981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5908_ _2829_ vssd1 vssd1 vccd1 vccd1 _2830_ sky130_fd_sc_hd__buf_4
X_6888_ clknet_leaf_83_core_clock _0149_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5839_ _2786_ vssd1 vssd1 vccd1 vccd1 _2787_ sky130_fd_sc_hd__buf_4
XANTENNA__6403__B _3118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7113__CLK clknet_leaf_33_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5734__S _2720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6479__A1 _1989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_3_core_clock_A clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_150_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3388__S1 _0864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input152_A c1_o_mem_high_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4874__A _2204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_78_core_clock_A clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input13_A c0_o_mem_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5206__A2 _2409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6313__B _3059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5390__A1 _2517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3953__A _1466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7425__A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3379__S1 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output636_A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4170_ _1676_ _1677_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__and2b_1
XFILLER_228_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4784__A _2150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3456__A1 _0918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput390 inner_wb_i_dat[10] vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_8
XFILLER_243_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3551__S1 _0902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6811_ clknet_leaf_85_core_clock _0072_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[14\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7136__CLK clknet_leaf_13_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6742_ clknet_leaf_67_core_clock _0003_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3954_ net313 _1416_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__nand2_1
XFILLER_223_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4950__C _2259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6673_ clknet_leaf_58_core_clock _0743_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6223__B _2118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_80_core_clock_A clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3885_ net254 _1401_ _1386_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__mux2_4
XANTENNA__3339__S _0865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4708__A1 _2016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5624_ _2240_ _2650_ _2660_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__a21o_1
XANTENNA__4024__A _1416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7286__CLK clknet_leaf_26_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5555_ _2242_ _2623_ _2625_ immu_0.page_table\[1\]\[7\] vssd1 vssd1 vccd1 vccd1 _0183_
+ sky130_fd_sc_hd__o22a_1
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4506_ _1979_ _1970_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__and2_1
XFILLER_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5486_ net93 _2577_ vssd1 vssd1 vccd1 vccd1 _2587_ sky130_fd_sc_hd__and2_1
XANTENNA__5133__A1 _2224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7225_ clknet_leaf_17_core_clock _0486_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4437_ _1926_ _1923_ vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__nor2_1
XFILLER_132_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7156_ clknet_leaf_29_core_clock _0417_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[9\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_258_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4368_ _1496_ _1869_ _1871_ _1530_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__o211a_1
XANTENNA__3695__A1 _0872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input5_A c0_o_instr_long_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6107_ _2799_ _2944_ vssd1 vssd1 vccd1 vccd1 _2951_ sky130_fd_sc_hd__and2_1
X_3319_ _0901_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__clkbuf_8
XFILLER_58_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7087_ clknet_leaf_93_core_clock _0348_ vssd1 vssd1 vccd1 vccd1 dmmu0.long_off_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_2_3_0_core_clock_A clknet_1_1_1_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4299_ _1413_ _1790_ _1794_ _1803_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__o31a_1
X_6038_ _2797_ _2904_ vssd1 vssd1 vccd1 vccd1 _2909_ sky130_fd_sc_hd__and2_1
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3447__B2 _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5302__B _2367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6414__A _1958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4947__A1 _1974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6133__B dmmu0.page_table\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3249__S _0847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6164__A3 _2981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5972__B _2861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3773__A _1336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6653__CLK clknet_leaf_39_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input367_A ic1_wb_adr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3712__S net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3438__A1 _0881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7159__CLK clknet_leaf_12_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3948__A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6324__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3670_ _1250_ _1251_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__nor2_1
XFILLER_118_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3683__A _0869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5340_ _2489_ immu_0.page_table\[9\]\[4\] _2495_ _2501_ vssd1 vssd1 vccd1 vccd1 _0092_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__3913__A2 _1426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5115__A1 _2347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5271_ _2217_ _2318_ vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_37_core_clock clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_181_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7010_ clknet_leaf_78_core_clock _0271_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4222_ _1413_ _1715_ _1719_ _1728_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__o31a_1
XANTENNA__4469__A3 _1924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4153_ _1454_ _1660_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__or2_1
XFILLER_256_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4084_ _1590_ _1592_ _1593_ _1530_ _1553_ vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__a221oi_2
XFILLER_283_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3429__B2 _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6526__CLK clknet_leaf_30_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6234__A _2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4680__C _2086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4986_ _2105_ vssd1 vssd1 vccd1 vccd1 _2284_ sky130_fd_sc_hd__buf_2
XFILLER_211_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6394__A3 _3116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3937_ _1450_ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__clkbuf_4
X_6725_ clknet_leaf_62_core_clock _0795_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[14\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinterconnect_inner_715 vssd1 vssd1 vccd1 vccd1 interconnect_inner_715/HI c0_i_core_int_sreg[6]
+ sky130_fd_sc_hd__conb_1
XANTENNA__3601__A1 _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinterconnect_inner_726 vssd1 vssd1 vccd1 vccd1 interconnect_inner_726/HI c1_i_core_int_sreg[3]
+ sky130_fd_sc_hd__conb_1
Xinterconnect_inner_737 vssd1 vssd1 vccd1 vccd1 interconnect_inner_737/HI c1_i_core_int_sreg[14]
+ sky130_fd_sc_hd__conb_1
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6656_ clknet_leaf_40_core_clock _0726_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_76_core_clock clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_core_clock
+ sky130_fd_sc_hd__clkbuf_16
X_3868_ _0812_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__buf_4
XFILLER_164_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5607_ _2649_ vssd1 vssd1 vccd1 vccd1 _2650_ sky130_fd_sc_hd__clkbuf_4
X_6587_ clknet_leaf_45_core_clock _0657_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4689__A _2000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3799_ net228 _1348_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__and2_1
XFILLER_191_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5538_ _2561_ vssd1 vssd1 vccd1 vccd1 _2618_ sky130_fd_sc_hd__buf_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5469_ _2576_ immu_0.page_table\[4\]\[1\] _2574_ _2578_ vssd1 vssd1 vccd1 vccd1 _0144_
+ sky130_fd_sc_hd__a31o_1
XFILLER_274_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput650 net650 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[12] sky130_fd_sc_hd__buf_2
Xoutput661 net661 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[8] sky130_fd_sc_hd__buf_2
Xoutput672 net672 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[16] sky130_fd_sc_hd__buf_2
XFILLER_278_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7208_ clknet_leaf_27_core_clock _0469_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[6\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5657__A2 _2669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput683 net683 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[4] sky130_fd_sc_hd__buf_2
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput694 net694 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[13] sky130_fd_sc_hd__buf_2
XFILLER_278_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7139_ clknet_leaf_33_core_clock _0400_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[10\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7301__CLK clknet_leaf_44_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4855__C _2197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5313__A _1937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5967__B _2861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input115_A c1_o_instr_long_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4363__S _1524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6144__A _2971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5593__A1 _2240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 c0_o_mem_addr[14] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_2
XFILLER_10_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input80_A c0_sr_bus_addr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput29 c0_o_mem_data[0] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_167_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5345__A1 _2503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4599__A _2038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5896__A2 _2812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6549__CLK clknet_leaf_48_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6038__B _2904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4084__B2 _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6699__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5596__C _2634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4840_ _1974_ _2189_ _2192_ immu_1.page_table\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 _0710_
+ sky130_fd_sc_hd__o22a_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _2150_ immu_1.page_table\[5\]\[9\] _2140_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__and3_1
XFILLER_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5584__A1 _2227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5893__A _2819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6510_ clknet_leaf_60_core_clock _0580_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3722_ _1256_ _1301_ _1300_ _0879_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__a31o_1
X_7490_ net180 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_1
XFILLER_173_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6441_ net199 _3136_ vssd1 vssd1 vccd1 vccd1 _3149_ sky130_fd_sc_hd__and2_1
XANTENNA__5336__A1 _2489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4139__A2 _1642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3653_ dmmu0.page_table\[4\]\[11\] dmmu0.page_table\[5\]\[11\] _0895_ vssd1 vssd1
+ vccd1 vccd1 _1235_ sky130_fd_sc_hd__mux2_1
XFILLER_173_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5887__A2 _2812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6372_ _3101_ dmmu1.page_table\[2\]\[8\] _3096_ _3108_ vssd1 vssd1 vccd1 vccd1 _0517_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__4302__A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3584_ _0893_ _1153_ _1162_ _1167_ _0879_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__o32a_2
XANTENNA__5117__B _2355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5323_ _2489_ immu_0.page_table\[10\]\[8\] _2480_ _2491_ vssd1 vssd1 vccd1 vccd1
+ _0085_ sky130_fd_sc_hd__a31o_1
XFILLER_114_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5254_ _2447_ dmmu0.page_table\[7\]\[5\] _2445_ vssd1 vssd1 vccd1 vccd1 _2452_ sky130_fd_sc_hd__and3_1
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4205_ immu_0.page_table\[4\]\[7\] immu_0.page_table\[5\]\[7\] _1472_ vssd1 vssd1
+ vccd1 vccd1 _1712_ sky130_fd_sc_hd__mux2_1
XFILLER_87_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5185_ _2400_ dmmu0.page_table\[9\]\[11\] _2391_ vssd1 vssd1 vccd1 vccd1 _2405_ sky130_fd_sc_hd__and3_1
XANTENNA__6229__A _2793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4136_ _1478_ _1643_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__or2_1
XFILLER_256_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4067_ net5 immu_0.high_addr_off\[0\] net2 vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__o21ai_1
XFILLER_283_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4691__B _2099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4969_ _1967_ _2274_ _2277_ immu_1.page_table\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 _0754_
+ sky130_fd_sc_hd__o22a_1
XFILLER_196_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6708_ clknet_leaf_61_core_clock _0778_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5327__A1 _2489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6639_ clknet_leaf_56_core_clock _0709_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3433__S0 _0858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput480 net480 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[5] sky130_fd_sc_hd__buf_2
Xoutput491 net491 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[14] sky130_fd_sc_hd__buf_2
XANTENNA__4838__B1 _2192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_17_core_clock_A clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4358__S _1439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6139__A _2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input232_A dcache_wb_adr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5978__A _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4882__A _2215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6841__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5802__A2 _2747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5566__A1 _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6991__CLK clknet_leaf_9_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5318__A1 _2363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3329__B1 _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3424__S0 _0897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output451_A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3975__S1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7433__A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4776__B _2153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3727__S1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6049__A _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5888__A _2681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6483__S _3172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4792__A _2150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6990_ clknet_leaf_8_core_clock _0251_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_253_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5941_ _2849_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_225_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5400__B _2527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5872_ _1991_ _2788_ vssd1 vssd1 vccd1 vccd1 _2809_ sky130_fd_sc_hd__and2_1
XFILLER_230_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3201__A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4823_ _2182_ immu_1.page_table\[2\]\[7\] _2174_ vssd1 vssd1 vccd1 vccd1 _2183_ sky130_fd_sc_hd__and3_1
XANTENNA__5557__A1 _1948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3568__B1 _0854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5021__A3 _2298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4754_ _2134_ immu_1.page_table\[5\]\[1\] _2140_ vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__and3_1
XFILLER_239_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3705_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__inv_2
X_7473_ net164 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_1
X_4685_ _2023_ _2083_ _2097_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__a21o_1
XANTENNA__6231__B _3021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3347__S _0858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5128__A _2216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3636_ dmmu0.page_table\[4\]\[10\] dmmu0.page_table\[5\]\[10\] dmmu0.page_table\[6\]\[10\]
+ dmmu0.page_table\[7\]\[10\] net15 net16 vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__mux4_1
X_6424_ _3128_ dmmu1.page_table\[0\]\[2\] _3135_ _3140_ vssd1 vssd1 vccd1 vccd1 _0537_
+ sky130_fd_sc_hd__a31o_1
XFILLER_174_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6714__CLK clknet_leaf_62_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6355_ _3085_ dmmu1.page_table\[2\]\[0\] _3096_ _3099_ vssd1 vssd1 vccd1 vccd1 _0509_
+ sky130_fd_sc_hd__a31o_1
XFILLER_127_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3567_ dmmu1.page_table\[10\]\[9\] dmmu1.page_table\[11\]\[9\] _1146_ vssd1 vssd1
+ vccd1 vccd1 _1151_ sky130_fd_sc_hd__mux2_1
XANTENNA__3871__A _1392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5306_ _1930_ _2367_ vssd1 vssd1 vccd1 vccd1 _2482_ sky130_fd_sc_hd__nor2_4
X_6286_ _3056_ vssd1 vssd1 vccd1 vccd1 _3057_ sky130_fd_sc_hd__clkbuf_2
XFILLER_88_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3498_ dmmu1.page_table\[8\]\[7\] dmmu1.page_table\[9\]\[7\] dmmu1.page_table\[10\]\[7\]
+ dmmu1.page_table\[11\]\[7\] _0891_ _0860_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__mux4_1
XFILLER_88_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_8_core_clock_A clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_248_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput208 c1_sr_bus_data_o[8] vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
X_5237_ _1912_ _2439_ vssd1 vssd1 vccd1 vccd1 _2440_ sky130_fd_sc_hd__or2_4
Xinput219 dcache_mem_o_data[14] vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_4
XANTENNA__6864__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5168_ _2384_ dmmu0.page_table\[9\]\[3\] _2392_ vssd1 vssd1 vccd1 vccd1 _2396_ sky130_fd_sc_hd__and3_1
XFILLER_271_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5798__A _2681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4119_ immu_1.page_table\[2\]\[5\] immu_1.page_table\[3\]\[5\] _1448_ vssd1 vssd1
+ vccd1 vccd1 _1628_ sky130_fd_sc_hd__mux2_1
XFILLER_17_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5099_ _1926_ _2352_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__nor2_1
XANTENNA__4048__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6406__B _3118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4207__A _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5548__A1 _2210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5012__A3 _2298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4220__A1 _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3257__S _0847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input182_A c1_sr_bus_addr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5980__B _2861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4877__A _2210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5720__A1 _2253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input43_A c0_o_mem_data[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5079__A3 _2336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4039__A1 _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5501__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4134__S1 _1570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5787__A1 _2232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7428__A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6332__A _2931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6737__CLK clknet_leaf_66_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_85_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_156_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4470_ net93 vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__buf_4
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3421_ net53 _1008_ _1009_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__a21o_1
X_6140_ _2239_ _2960_ _2969_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__a21o_1
XFILLER_143_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ _0864_ _0943_ _0880_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__mux2_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6071_ _2797_ _2924_ vssd1 vssd1 vccd1 vccd1 _2929_ sky130_fd_sc_hd__and2_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ net155 net154 net157 net156 vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__or4_1
XFILLER_97_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _1937_ _2302_ vssd1 vssd1 vccd1 vccd1 _2306_ sky130_fd_sc_hd__and2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3630__S net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5411__A _1930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6973_ clknet_leaf_0_core_clock _0234_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[11\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_213_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5924_ _2834_ dmmu0.page_table\[5\]\[6\] _2832_ vssd1 vssd1 vccd1 vccd1 _2840_ sky130_fd_sc_hd__and3_1
XFILLER_241_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4450__A1 _1911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5855_ _2618_ dmmu1.page_table\[15\]\[4\] _2787_ _2798_ vssd1 vssd1 vccd1 vccd1 _0310_
+ sky130_fd_sc_hd__a31o_1
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6242__A _2891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4806_ _2084_ _2170_ vssd1 vssd1 vccd1 vccd1 _2173_ sky130_fd_sc_hd__or2_1
XANTENNA__5784__C _2751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5786_ _2749_ dmmu0.page_table\[13\]\[4\] _2751_ vssd1 vssd1 vccd1 vccd1 _2756_ sky130_fd_sc_hd__and3_1
XANTENNA__3636__S0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5950__A1 _1940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4737_ _2016_ _2120_ _2130_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__a21o_1
XANTENNA__4753__A2 _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4668_ _2006_ _2083_ _2088_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__a21o_1
X_7456_ net389 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3619_ _0868_ _1201_ net122 vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__o21a_1
X_6407_ _3128_ dmmu1.page_table\[1\]\[9\] _3116_ _3129_ vssd1 vssd1 vccd1 vccd1 _0531_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__4697__A _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4599_ _2038_ immu_1.page_table\[13\]\[10\] _2031_ vssd1 vssd1 vccd1 vccd1 _2044_
+ sky130_fd_sc_hd__and3_1
XFILLER_134_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7387_ net357 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4061__S0 _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6338_ _3085_ dmmu1.page_table\[3\]\[7\] _3077_ _3088_ vssd1 vssd1 vccd1 vccd1 _0503_
+ sky130_fd_sc_hd__a31o_1
XFILLER_103_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6269_ _3042_ dmmu1.page_table\[5\]\[5\] _3038_ _3047_ vssd1 vssd1 vccd1 vccd1 _0475_
+ sky130_fd_sc_hd__a31o_1
XFILLER_76_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5481__A3 _2574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6417__A _2784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4863__C _2197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7192__CLK clknet_leaf_27_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4992__A2 _2280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5694__C _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6152__A _2971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6194__A1 _2994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input397_A inner_wb_i_dat[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5991__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3952__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6046__B _2904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3970_ _1478_ _1482_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__nand2_1
XFILLER_250_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6185__A1 _2994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5640_ _1914_ _2215_ vssd1 vssd1 vccd1 vccd1 _2670_ sky130_fd_sc_hd__or2_2
XFILLER_203_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5571_ _2242_ _2627_ _2630_ immu_0.page_table\[0\]\[7\] vssd1 vssd1 vccd1 vccd1 _0194_
+ sky130_fd_sc_hd__o22a_1
XFILLER_176_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4735__A2 _2120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4522_ _1976_ dmmu1.page_table\[14\]\[10\] _1963_ _1990_ vssd1 vssd1 vccd1 vccd1
+ _0594_ sky130_fd_sc_hd__a31o_1
XFILLER_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7310_ clknet_leaf_3_core_clock _0571_ vssd1 vssd1 vccd1 vccd1 dmmu1.long_off_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7241_ clknet_leaf_24_core_clock _0502_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4453_ _1911_ immu_0.page_table\[11\]\[4\] _1924_ _1938_ vssd1 vssd1 vccd1 vccd1
+ _0577_ sky130_fd_sc_hd__a31o_1
XFILLER_236_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4043__S0 _1453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4948__C _2259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3404_ _0839_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__clkbuf_4
XFILLER_104_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7172_ clknet_leaf_37_core_clock _0433_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4384_ _1831_ _1835_ _1886_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__a21o_1
XANTENNA__7065__CLK clknet_leaf_11_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6123_ _2216_ _2621_ vssd1 vssd1 vccd1 vccd1 _2959_ sky130_fd_sc_hd__nor2_1
X_3335_ net1 net53 vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__nor2_2
XFILLER_124_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6054_ _2914_ dmmu1.page_table\[11\]\[11\] _2901_ _2917_ vssd1 vssd1 vccd1 vccd1
+ _0390_ sky130_fd_sc_hd__a31o_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ net121 vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__clkbuf_4
XFILLER_218_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _2284_ immu_1.page_table\[15\]\[10\] _2281_ vssd1 vssd1 vccd1 vccd1 _2294_
+ sky130_fd_sc_hd__and3_1
XANTENNA__4120__B1 _1451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3197_ mem_dcache_arb.select net562 _0817_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__o21a_2
XFILLER_54_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4671__A1 _2008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6902__CLK clknet_leaf_79_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4980__A _1999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6956_ clknet_leaf_85_core_clock _0217_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5907_ _2216_ _2555_ vssd1 vssd1 vccd1 vccd1 _2829_ sky130_fd_sc_hd__nor2_2
XANTENNA__4974__A2 _2274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6887_ clknet_leaf_84_core_clock _0148_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3596__A _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6176__A1 _2977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5838_ _2785_ vssd1 vssd1 vccd1 vccd1 _2786_ sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5923__A1 _2235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5769_ _2736_ dmmu0.page_table\[4\]\[11\] _2731_ vssd1 vssd1 vccd1 vccd1 _2745_ sky130_fd_sc_hd__and3_1
XFILLER_194_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7508_ net395 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7439_ net68 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_1
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input145_A c1_o_mem_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4366__S _1438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5454__A3 _2557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4593__C _2032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5051__A _1935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input312_A ic0_wb_adr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6582__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5986__A _1993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4890__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7088__CLK clknet_leaf_2_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_core_clock clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4025__S0 _1472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5678__A0 _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4768__C _2140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4130__A _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output531_A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output629_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7441__A net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6057__A _1958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput380 ic1_wb_sel[0] vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_1
Xinput391 inner_wb_i_dat[11] vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_6
XFILLER_282_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6810_ clknet_leaf_87_core_clock _0071_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6491__S _3172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6741_ clknet_leaf_66_core_clock _0002_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3953_ _1466_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6672_ clknet_leaf_58_core_clock _0742_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3884_ net324 net378 _1390_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__mux2_1
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_66_core_clock clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4708__A2 _2101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5623_ _2655_ dmmu0.page_table\[15\]\[6\] _2652_ vssd1 vssd1 vccd1 vccd1 _2660_ sky130_fd_sc_hd__and3_1
X_5554_ _2239_ _2623_ _2625_ immu_0.page_table\[1\]\[6\] vssd1 vssd1 vccd1 vccd1 _0182_
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4505_ net205 vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__buf_6
X_5485_ _2576_ immu_0.page_table\[4\]\[9\] _2574_ _2586_ vssd1 vssd1 vccd1 vccd1 _0152_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__3355__S _0918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4678__C _2086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5136__A _2371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4436_ _1925_ vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__buf_4
XFILLER_144_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7224_ clknet_leaf_17_core_clock _0485_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5133__A2 _2369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7155_ clknet_leaf_30_core_clock _0416_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[9\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_4367_ _1584_ _1870_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__or2_1
XFILLER_98_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6106_ _2948_ dmmu1.page_table\[9\]\[4\] _2942_ _2950_ vssd1 vssd1 vccd1 vccd1 _0409_
+ sky130_fd_sc_hd__a31o_1
X_3318_ dmmu0.page_table\[14\]\[0\] dmmu0.page_table\[15\]\[0\] _0910_ vssd1 vssd1
+ vccd1 vccd1 _0911_ sky130_fd_sc_hd__mux2_1
X_7086_ clknet_leaf_0_core_clock _0347_ vssd1 vssd1 vccd1 vccd1 dmmu0.long_off_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4298_ _1535_ _1796_ _1798_ _1434_ _1802_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__a311o_1
XFILLER_112_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4186__S _1443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3249_ net129 net24 _0847_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__mux2_2
X_6037_ _2898_ dmmu1.page_table\[11\]\[3\] _2902_ _2908_ vssd1 vssd1 vccd1 vccd1 _0382_
+ sky130_fd_sc_hd__a31o_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4644__A1 _2010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6939_ clknet_leaf_82_core_clock _0200_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4947__A2 _2257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6414__B _2272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6149__A1 _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4215__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6133__C _2962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5046__A _1930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input262_A dcache_wb_o_dat[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6948__CLK clknet_leaf_81_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6388__A1 _3112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3948__B net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6324__B _3079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5060__A1 _2316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_24_core_clock_A clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_158_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output481_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7436__A net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5882__C _2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4020__C1 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5270_ _2253_ _2441_ _2460_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__a21o_1
XFILLER_141_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6312__A1 _3069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4221_ _1434_ _1723_ _1727_ _1410_ vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__o31a_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3903__S _1416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4152_ immu_1.page_table\[8\]\[6\] immu_1.page_table\[9\]\[6\] _1437_ vssd1 vssd1
+ vccd1 vccd1 _1660_ sky130_fd_sc_hd__mux2_1
XFILLER_256_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5418__A3 _2541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7103__CLK clknet_leaf_30_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4083_ immu_1.page_table\[0\]\[4\] immu_1.page_table\[1\]\[4\] immu_1.page_table\[2\]\[4\]
+ immu_1.page_table\[3\]\[4\] _1439_ _1496_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__mux4_1
XFILLER_228_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4626__A1 _2023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3204__A _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6234__B _3021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4985_ _1995_ _2280_ _2283_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__a21o_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6724_ clknet_leaf_61_core_clock _0794_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[14\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3936_ net368 vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__inv_2
Xinterconnect_inner_716 vssd1 vssd1 vccd1 vccd1 interconnect_inner_716/HI c0_i_core_int_sreg[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_176_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinterconnect_inner_727 vssd1 vssd1 vccd1 vccd1 interconnect_inner_727/HI c1_i_core_int_sreg[4]
+ sky130_fd_sc_hd__conb_1
Xinterconnect_inner_738 vssd1 vssd1 vccd1 vccd1 interconnect_inner_738/HI c1_i_core_int_sreg[15]
+ sky130_fd_sc_hd__conb_1
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6655_ clknet_leaf_39_core_clock _0725_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3867_ _1389_ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_1
XFILLER_149_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3874__A _1394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6250__A _1993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5792__C _2751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5606_ _2217_ _2296_ vssd1 vssd1 vccd1 vccd1 _2649_ sky130_fd_sc_hd__nor2_1
XFILLER_258_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6586_ clknet_leaf_45_core_clock _0656_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4689__B _2099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3798_ _1350_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_1
XFILLER_164_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5537_ _2603_ immu_0.page_table\[2\]\[8\] _2607_ _2617_ vssd1 vssd1 vccd1 vccd1 _0173_
+ sky130_fd_sc_hd__a31o_1
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6303__A1 _3053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput640 net640 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[9] sky130_fd_sc_hd__buf_2
X_5468_ net96 _2577_ vssd1 vssd1 vccd1 vccd1 _2578_ sky130_fd_sc_hd__and2_1
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput651 net651 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[13] sky130_fd_sc_hd__buf_2
XFILLER_2_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7207_ clknet_leaf_27_core_clock _0468_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[6\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_274_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput662 net662 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[9] sky130_fd_sc_hd__buf_2
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput673 net673 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[17] sky130_fd_sc_hd__buf_2
X_4419_ _1909_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_1
Xoutput684 net684 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[5] sky130_fd_sc_hd__buf_2
Xoutput695 net695 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[14] sky130_fd_sc_hd__buf_2
XFILLER_259_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5399_ _2531_ immu_0.page_table\[7\]\[7\] _2525_ _2535_ vssd1 vssd1 vccd1 vccd1 _0117_
+ sky130_fd_sc_hd__a31o_1
XFILLER_160_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7138_ clknet_leaf_28_core_clock _0399_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_246_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5313__B _2482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4078__C1 _1457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7069_ clknet_leaf_4_core_clock _0330_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[6\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6082__A3 _2922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5290__A1 _2243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input108_A c1_o_c_instr_page vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6620__CLK clknet_leaf_53_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5593__A2 _2632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3784__A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput19 c0_o_mem_addr[15] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_167_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6160__A _2982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input73_A c0_o_req_addr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5207__C _2411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7126__CLK clknet_leaf_33_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3723__S _0857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4856__A1 _1967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7276__CLK clknet_leaf_22_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3959__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6335__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5584__A2 _2632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4770_ _2105_ vssd1 vssd1 vccd1 vccd1 _2150_ sky130_fd_sc_hd__buf_2
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3721_ _1256_ _1300_ _1301_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__a21oi_1
XFILLER_186_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6440_ _1898_ dmmu1.page_table\[0\]\[10\] _3134_ _3148_ vssd1 vssd1 vccd1 vccd1 _0545_
+ sky130_fd_sc_hd__a31o_1
XFILLER_186_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3652_ dmmu0.page_table\[6\]\[11\] dmmu0.page_table\[7\]\[11\] _0896_ vssd1 vssd1
+ vccd1 vccd1 _1234_ sky130_fd_sc_hd__mux2_1
XFILLER_146_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6371_ net208 _3098_ vssd1 vssd1 vccd1 vccd1 _3108_ sky130_fd_sc_hd__and2_1
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3583_ _1165_ _1166_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5322_ _2310_ _2482_ vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__and2_1
XFILLER_173_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5253_ _2233_ _2442_ _2451_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__a21o_1
XANTENNA__4847__A1 _1989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4956__C _2259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5414__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4204_ _1707_ _1708_ _1709_ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__nand3_1
X_5184_ _2249_ _2389_ _2404_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__a21o_1
XANTENNA__6229__B _3021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4135_ immu_0.page_table\[2\]\[6\] immu_0.page_table\[3\]\[6\] _1601_ vssd1 vssd1
+ vccd1 vccd1 _1643_ sky130_fd_sc_hd__mux2_1
XFILLER_56_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_92_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__6064__A3 _2922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4066_ net5 immu_0.high_addr_off\[0\] vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__and2_1
XFILLER_271_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6643__CLK clknet_leaf_39_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4968_ _2275_ vssd1 vssd1 vccd1 vccd1 _2277_ sky130_fd_sc_hd__buf_4
XANTENNA__4378__A3 _1880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6793__CLK clknet_leaf_80_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6707_ clknet_leaf_62_core_clock _0777_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3919_ _1430_ _1431_ _1432_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__a21oi_1
X_4899_ _2229_ vssd1 vssd1 vccd1 vccd1 _2230_ sky130_fd_sc_hd__buf_4
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6638_ clknet_leaf_42_core_clock _0708_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3338__A1 _0890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3338__B2 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6569_ clknet_leaf_49_core_clock _0639_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[11\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_285_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3433__S1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput470 net470 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[10] sky130_fd_sc_hd__buf_2
XANTENNA__4838__A1 _1967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput481 net481 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[6] sky130_fd_sc_hd__buf_2
XANTENNA__4866__C _2197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5324__A _2312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput492 net492 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[15] sky130_fd_sc_hd__buf_2
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7299__CLK clknet_leaf_44_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5978__B _2861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input225_A dcache_mem_o_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5263__A1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3779__A _1340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6155__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5994__A _2879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4223__C1 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3577__A1 _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4403__A _1901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3329__A1 _0918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5869__A3 _2787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3424__S1 _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6516__CLK clknet_leaf_36_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output444_A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6049__B _2904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3501__A1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6065__A _2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5940_ dmmu0.long_off_reg\[0\] net92 _2848_ vssd1 vssd1 vccd1 vccd1 _2849_ sky130_fd_sc_hd__mux2_1
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5871_ _2805_ dmmu1.page_table\[15\]\[10\] _2786_ _2808_ vssd1 vssd1 vccd1 vccd1
+ _0316_ sky130_fd_sc_hd__a31o_1
XFILLER_33_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5006__A1 _1989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3201__B _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4822_ _2105_ vssd1 vssd1 vccd1 vccd1 _2182_ sky130_fd_sc_hd__buf_2
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5557__A2 _2623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3568__A1 _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4753_ _1996_ _2138_ _2141_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__a21o_1
XFILLER_159_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5409__A _1925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3704_ dmmu0.page_table\[8\]\[12\] dmmu0.page_table\[9\]\[12\] dmmu0.page_table\[10\]\[12\]
+ dmmu0.page_table\[11\]\[12\] net15 net16 vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__mux4_1
X_7472_ clknet_opt_2_1_core_clock vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__buf_2
X_4684_ _2089_ immu_1.page_table\[10\]\[9\] _2086_ vssd1 vssd1 vccd1 vccd1 _2097_
+ sky130_fd_sc_hd__and3_1
XANTENNA__5128__B _2367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6423_ net202 _3137_ vssd1 vssd1 vccd1 vccd1 _3140_ sky130_fd_sc_hd__and2_1
X_3635_ dmmu0.page_table\[0\]\[10\] dmmu0.page_table\[1\]\[10\] dmmu0.page_table\[2\]\[10\]
+ dmmu0.page_table\[3\]\[10\] _0895_ net16 vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__mux4_1
XFILLER_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6354_ net197 _3098_ vssd1 vssd1 vccd1 vccd1 _3099_ sky130_fd_sc_hd__and2_1
X_3566_ _0868_ _1149_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__and2_1
X_5305_ _2363_ immu_0.page_table\[10\]\[0\] _2480_ _2481_ vssd1 vssd1 vccd1 vccd1
+ _0077_ sky130_fd_sc_hd__a31o_1
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6285_ _2919_ _2153_ vssd1 vssd1 vccd1 vccd1 _3056_ sky130_fd_sc_hd__or2_1
X_3497_ dmmu1.page_table\[12\]\[7\] dmmu1.page_table\[13\]\[7\] dmmu1.page_table\[14\]\[7\]
+ dmmu1.page_table\[15\]\[7\] _0891_ _0860_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__mux4_1
XANTENNA__5144__A _2371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput209 c1_sr_bus_data_o[9] vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_4
X_5236_ net85 net84 vssd1 vssd1 vccd1 vccd1 _2439_ sky130_fd_sc_hd__or2b_1
XANTENNA__5493__A1 _2588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5167_ _2227_ _2390_ _2395_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__a21o_1
XFILLER_68_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4118_ _1442_ _1626_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__or2_1
XANTENNA__6037__A3 _2902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5098_ _2352_ vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__clkbuf_4
XFILLER_284_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4194__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4049_ immu_1.page_table\[14\]\[3\] immu_1.page_table\[15\]\[3\] _1493_ vssd1 vssd1
+ vccd1 vccd1 _1560_ sky130_fd_sc_hd__mux2_1
XFILLER_71_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5548__A2 _2623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3559__A1 _1088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5319__A _2300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6539__CLK clknet_leaf_48_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6141__C _2962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input175_A c1_o_req_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6689__CLK clknet_leaf_39_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3273__S _0865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input342_A ic1_mem_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input36_A c0_o_mem_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4039__A2 _1547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5501__B _2593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5787__A2 _2748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3302__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6200__A3 _3000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3448__S _0898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5229__A _2099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output561_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7444__A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3420_ net53 net1 vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__and2b_1
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3351_ _0934_ _0936_ _0938_ _0942_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__o22a_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6267__A3 _3038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3282_ _0855_ _0862_ _0867_ _0873_ _0874_ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__a221o_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6070_ _2914_ dmmu1.page_table\[10\]\[3\] _2922_ _2928_ vssd1 vssd1 vccd1 vccd1 _0395_
+ sky130_fd_sc_hd__a31o_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5475__A1 _2576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5899__A _2819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _2301_ immu_0.page_table\[15\]\[3\] _2298_ _2305_ vssd1 vssd1 vccd1 vccd1
+ _0778_ sky130_fd_sc_hd__a31o_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6019__A3 _2877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5227__A1 _2210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5411__B _2539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3238__A0 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4308__A _1584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6972_ clknet_leaf_88_core_clock _0233_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[11\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_253_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3212__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5130__C _2373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5923_ _2235_ _2830_ _2839_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__a21o_1
XFILLER_241_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5854_ _2797_ _2789_ vssd1 vssd1 vccd1 vccd1 _2798_ sky130_fd_sc_hd__and2_1
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4805_ _2171_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__6242__B _3021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5785_ _2229_ _2748_ _2755_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__a21o_1
XFILLER_21_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3358__S _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3636__S1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4736_ _2121_ immu_1.page_table\[6\]\[6\] _2123_ vssd1 vssd1 vccd1 vccd1 _2130_ sky130_fd_sc_hd__and3_1
XFILLER_174_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7455_ net710 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_1
XFILLER_119_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4667_ _2072_ immu_1.page_table\[10\]\[1\] _2086_ vssd1 vssd1 vccd1 vccd1 _2088_
+ sky130_fd_sc_hd__and3_1
XFILLER_119_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6406_ net209 _3118_ vssd1 vssd1 vccd1 vccd1 _3129_ sky130_fd_sc_hd__and2_1
XANTENNA__6831__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3618_ dmmu1.page_table\[14\]\[10\] dmmu1.page_table\[15\]\[10\] net120 vssd1 vssd1
+ vccd1 vccd1 _1201_ sky130_fd_sc_hd__mux2_1
X_7386_ net356 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_1
X_4598_ _2023_ _2030_ _2043_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__a21o_1
XANTENNA__4061__S1 _1570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4189__S _1443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6337_ net207 _3079_ vssd1 vssd1 vccd1 vccd1 _3088_ sky130_fd_sc_hd__and2_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3549_ _1132_ _1133_ _0957_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__o21ai_1
XFILLER_249_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6258__A3 _3038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6268_ _2799_ _3040_ vssd1 vssd1 vccd1 vccd1 _3047_ sky130_fd_sc_hd__and2_1
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5219_ _2416_ dmmu0.page_table\[8\]\[12\] _2410_ vssd1 vssd1 vccd1 vccd1 _2425_ sky130_fd_sc_hd__and3_1
XFILLER_229_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6199_ _2795_ _3002_ vssd1 vssd1 vccd1 vccd1 _3006_ sky130_fd_sc_hd__and2_1
XANTENNA__5602__A _2640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6417__B _2272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5218__A1 _2251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4977__B1 _2277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6430__A3 _3135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5049__A _1933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input292_A ic0_mem_data[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_core_clock_A clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_200_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4888__A _2204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3792__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_17_core_clock clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_153_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3704__A1 dmmu0.page_table\[9\]\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6249__A3 _3018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3731__S net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4128__A _1570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output407_A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6704__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_core_clock clknet_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_1_0_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_223_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3967__A _1472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7439__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6343__A _2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_56_core_clock clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4196__A1 _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6854__CLK clknet_leaf_70_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5570_ _2239_ _2627_ _2630_ immu_0.page_table\[0\]\[6\] vssd1 vssd1 vccd1 vccd1 _0193_
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4521_ _1989_ _1970_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__and2_1
XFILLER_144_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6489__S _3172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7240_ clknet_leaf_20_core_clock _0501_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4452_ _1937_ _1931_ vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__and2_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4043__S1 _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3403_ _0980_ _0984_ _0988_ _0992_ vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__o22a_4
X_7171_ clknet_leaf_33_core_clock _0432_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4383_ net12 immu_0.high_addr_off\[7\] vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__xor2_1
XANTENNA__3207__A _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6122_ _2948_ dmmu1.page_table\[9\]\[12\] _2941_ _2958_ vssd1 vssd1 vccd1 vccd1 _0417_
+ sky130_fd_sc_hd__a31o_1
X_3334_ net53 _0926_ vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__and2_1
XANTENNA__5448__A1 _2562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6053_ _1991_ _2903_ vssd1 vssd1 vccd1 vccd1 _2917_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_31_core_clock_A clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3265_ _0857_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__buf_6
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _1987_ _2280_ _2293_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__a21o_1
XANTENNA__4120__A1 _1584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3554__S0 _0896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3196_ mem_dcache_arb.transfer_active _0809_ _0816_ vssd1 vssd1 vccd1 vccd1 _0817_
+ sky130_fd_sc_hd__or3_2
XFILLER_273_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4671__A2 _2083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4980__B _2278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6955_ clknet_leaf_85_core_clock _0216_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_214_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3877__A _1396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5620__A1 _2233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5906_ net95 _2811_ _2828_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__a21o_1
XFILLER_241_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6886_ clknet_leaf_71_core_clock _0147_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3596__B _1179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5837_ _2784_ _2278_ vssd1 vssd1 vccd1 vccd1 _2785_ sky130_fd_sc_hd__or2_1
XFILLER_194_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5923__A2 _2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5768_ _1950_ _2729_ _2744_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__a21o_1
XFILLER_277_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7507_ net394 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_1
XFILLER_147_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4719_ _2000_ _2118_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__nor2_1
XFILLER_194_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5699_ _2227_ _2700_ _2705_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__a21o_1
XFILLER_30_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4501__A _1898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7438_ net67 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_1
XFILLER_107_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7369_ net293 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_2
XFILLER_162_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5332__A _1930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input138_A c1_o_mem_data[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6727__CLK clknet_leaf_66_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5051__B _2322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3870__A0 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input305_A ic0_mem_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5611__A1 _2211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6163__A _2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6877__CLK clknet_leaf_70_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5390__A3 _2525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5507__A net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4025__S1 _1419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output524_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3461__S _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4784__C _2157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput370 ic1_wb_adr[1] vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_1
XFILLER_208_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput381 ic1_wb_sel[1] vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_1
Xinput392 inner_wb_i_dat[12] vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_6
XFILLER_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3861__A0 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4292__S _1425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6740_ clknet_leaf_66_core_clock _0001_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6073__A _2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3952_ net234 _1465_ _0811_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__mux2_4
XFILLER_223_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6671_ clknet_leaf_4_core_clock _0741_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_3883_ _1400_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_1
XFILLER_188_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5622_ _2236_ _2650_ _2659_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__a21o_1
XFILLER_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7032__CLK clknet_leaf_13_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5553_ _2235_ _2623_ _2625_ immu_0.page_table\[1\]\[5\] vssd1 vssd1 vccd1 vccd1 _0181_
+ sky130_fd_sc_hd__o22a_1
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5417__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4504_ _1976_ dmmu1.page_table\[14\]\[4\] _1964_ _1978_ vssd1 vssd1 vccd1 vccd1 _0588_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__4321__A _1581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5484_ net104 _2577_ vssd1 vssd1 vccd1 vccd1 _2586_ sky130_fd_sc_hd__and2_1
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5669__A1 _2253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7223_ clknet_leaf_23_core_clock _0484_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4435_ net92 vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__inv_2
XFILLER_144_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7182__CLK clknet_leaf_29_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7154_ clknet_leaf_29_core_clock _0415_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[9\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_258_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4366_ immu_1.page_table\[2\]\[10\] immu_1.page_table\[3\]\[10\] _1438_ vssd1 vssd1
+ vccd1 vccd1 _1870_ sky130_fd_sc_hd__mux2_1
XFILLER_263_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6105_ _2797_ _2944_ vssd1 vssd1 vccd1 vccd1 _2950_ sky130_fd_sc_hd__and2_1
X_3317_ _0900_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__buf_6
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6248__A _1991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7085_ clknet_leaf_93_core_clock _0346_ vssd1 vssd1 vccd1 vccd1 dmmu0.long_off_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4297_ _1424_ _1799_ _1801_ _1432_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__o211a_1
XANTENNA__3371__S _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6036_ _2795_ _2904_ vssd1 vssd1 vccd1 vccd1 _2908_ sky130_fd_sc_hd__and2_1
X_3248_ _0839_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__buf_4
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4991__A _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6938_ clknet_leaf_84_core_clock _0199_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6869_ clknet_leaf_69_core_clock _0130_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[6\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_222_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5046__B _2318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input255_A dcache_wb_cyc vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6158__A _2980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4406__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7055__CLK clknet_leaf_30_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4125__B _1633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_core_clock clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_158_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4020__B1 _1528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4571__A1 _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4141__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5115__A3 _2353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3980__A _1443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7452__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4323__A1 _1457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4220_ _1423_ _1724_ _1726_ _1416_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__o211a_1
X_4151_ immu_1.page_table\[10\]\[6\] immu_1.page_table\[11\]\[6\] _1453_ vssd1 vssd1
+ vccd1 vccd1 _1659_ sky130_fd_sc_hd__mux2_1
XANTENNA__4287__S _1425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4082_ _1523_ _1591_ _1516_ vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__o21a_1
XFILLER_228_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4626__A2 _2047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5700__A _2682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4316__A _1584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4984_ _2262_ immu_1.page_table\[15\]\[0\] _2282_ vssd1 vssd1 vccd1 vccd1 _2283_
+ sky130_fd_sc_hd__and3_1
XFILLER_211_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3220__A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6723_ clknet_leaf_63_core_clock _0793_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3935_ immu_1.page_table\[4\]\[0\] immu_1.page_table\[5\]\[0\] _1448_ vssd1 vssd1
+ vccd1 vccd1 _1449_ sky130_fd_sc_hd__mux2_1
Xinterconnect_inner_717 vssd1 vssd1 vccd1 vccd1 interconnect_inner_717/HI c0_i_core_int_sreg[8]
+ sky130_fd_sc_hd__conb_1
Xinterconnect_inner_728 vssd1 vssd1 vccd1 vccd1 interconnect_inner_728/HI c1_i_core_int_sreg[5]
+ sky130_fd_sc_hd__conb_1
X_6654_ clknet_leaf_40_core_clock _0724_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xinterconnect_inner_739 vssd1 vssd1 vccd1 vccd1 interconnect_inner_739/HI c1_i_irq
+ sky130_fd_sc_hd__conb_1
X_3866_ net248 _1388_ _1386_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__mux2_4
XANTENNA__6000__A1 _2884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5605_ _2253_ _2631_ _2648_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__a21o_1
XFILLER_137_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6250__B _3020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6585_ clknet_leaf_46_core_clock _0655_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3797_ net227 _1348_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__and2_1
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4562__A1 _2019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4051__A _1442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5536_ net103 _2609_ vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__and2_1
XANTENNA__6572__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4986__A _2105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5467_ _1922_ _2572_ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__nor2_4
XFILLER_274_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput630 net630 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[14] sky130_fd_sc_hd__buf_2
XFILLER_132_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput641 net641 vssd1 vssd1 vccd1 vccd1 ic1_mem_cache_flush sky130_fd_sc_hd__buf_2
X_7206_ clknet_leaf_27_core_clock _0467_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[6\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_278_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput652 net652 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[14] sky130_fd_sc_hd__buf_2
Xoutput663 net663 vssd1 vssd1 vccd1 vccd1 inner_wb_4_burst sky130_fd_sc_hd__buf_2
X_4418_ _1373_ net230 vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__and2_4
Xoutput674 net674 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[18] sky130_fd_sc_hd__buf_2
X_5398_ _1944_ _2527_ vssd1 vssd1 vccd1 vccd1 _2535_ sky130_fd_sc_hd__and2_1
Xoutput685 net685 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[6] sky130_fd_sc_hd__buf_2
XFILLER_132_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput696 net696 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[15] sky130_fd_sc_hd__buf_2
XFILLER_207_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7137_ clknet_leaf_34_core_clock _0398_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4349_ _1432_ _1846_ _1848_ _1413_ _1852_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__a311o_1
XFILLER_247_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7068_ clknet_leaf_4_core_clock _0329_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[6\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5814__A1 _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6019_ _2884_ dmmu1.page_table\[12\]\[10\] _2877_ _2896_ vssd1 vssd1 vccd1 vccd1
+ _0376_ sky130_fd_sc_hd__a31o_1
XFILLER_100_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5610__A _2640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5290__A2 _2462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7078__CLK clknet_leaf_11_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6425__B _3137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4226__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6144__C _2962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6441__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3784__B _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6915__CLK clknet_leaf_76_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5345__A3 _2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5057__A _1942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input372_A ic1_wb_adr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input66_A c0_o_req_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4896__A _2204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4856__A2 _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3305__A _0897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6335__B _3079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4136__A _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6230__A1 _3010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7447__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3720_ net157 dmmu1.long_off_reg\[7\] vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__xor2_1
XANTENNA__5893__C _2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6595__CLK clknet_leaf_59_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3651_ _0908_ _1230_ _1232_ _0917_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__o211a_1
XFILLER_146_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5336__A3 _2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6370_ _3101_ dmmu1.page_table\[2\]\[7\] _3096_ _3107_ vssd1 vssd1 vccd1 vccd1 _0516_
+ sky130_fd_sc_hd__a31o_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3582_ _1124_ _1125_ _1123_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__a21bo_1
XFILLER_127_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5321_ _2489_ immu_0.page_table\[10\]\[7\] _2480_ _2490_ vssd1 vssd1 vccd1 vccd1
+ _0084_ sky130_fd_sc_hd__a31o_1
XFILLER_127_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6497__S _3172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3914__S _1408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6297__A1 _3053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5252_ _2447_ dmmu0.page_table\[7\]\[4\] _2445_ vssd1 vssd1 vccd1 vccd1 _2451_ sky130_fd_sc_hd__and3_1
XFILLER_244_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5414__B _2543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4203_ _1707_ _1708_ _1709_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__a21o_1
X_5183_ _2400_ dmmu0.page_table\[9\]\[10\] _2391_ vssd1 vssd1 vccd1 vccd1 _2404_ sky130_fd_sc_hd__and3_1
XFILLER_229_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4134_ immu_0.page_table\[4\]\[6\] immu_0.page_table\[5\]\[6\] immu_0.page_table\[6\]\[6\]
+ immu_0.page_table\[7\]\[6\] _1409_ _1570_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__mux4_2
XFILLER_110_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7220__CLK clknet_leaf_27_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4065_ _1571_ _1572_ _1573_ _1574_ _1479_ _1413_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__mux4_2
XFILLER_283_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4967_ _1965_ _2274_ _2276_ immu_1.page_table\[0\]\[0\] vssd1 vssd1 vccd1 vccd1 _0753_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_212_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3918_ net314 vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__clkbuf_4
X_6706_ clknet_leaf_61_core_clock _0776_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4783__A1 _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4898_ net98 vssd1 vssd1 vccd1 vccd1 _2229_ sky130_fd_sc_hd__buf_6
XFILLER_132_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6637_ clknet_leaf_57_core_clock _0707_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3849_ _1373_ net260 vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__and2_4
XFILLER_192_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3338__A2 _0894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6568_ clknet_leaf_49_core_clock _0638_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[11\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5519_ _1925_ _2606_ vssd1 vssd1 vccd1 vccd1 _2608_ sky130_fd_sc_hd__nor2_1
XFILLER_145_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6499_ _1914_ _1919_ _2426_ vssd1 vssd1 vccd1 vccd1 _3181_ sky130_fd_sc_hd__or3_1
XFILLER_279_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput460 net460 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[9] sky130_fd_sc_hd__buf_2
XFILLER_105_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput471 net471 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[11] sky130_fd_sc_hd__buf_2
XANTENNA__4838__A2 _2189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput482 net482 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[7] sky130_fd_sc_hd__buf_2
XANTENNA__5324__B _2482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput493 net493 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[16] sky130_fd_sc_hd__buf_2
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6139__C _2962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5263__A2 _2442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input120_A c1_o_mem_addr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6155__B net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input218_A dcache_mem_o_data[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5994__B _2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4223__B1 _1729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3795__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4774__A1 _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6171__A _2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5318__A3 _2480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3734__C1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6279__A1 _3042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output437_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_36_core_clock_A clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4792__C _2157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5250__A _2447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6065__B _2924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5870_ _1989_ _2788_ vssd1 vssd1 vccd1 vccd1 _2808_ sky130_fd_sc_hd__and2_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4821_ _2016_ _2172_ _2181_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__a21o_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6081__A _2891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4752_ _2134_ immu_1.page_table\[5\]\[0\] _2140_ vssd1 vssd1 vccd1 vccd1 _2141_ sky130_fd_sc_hd__and3_1
XANTENNA__4765__A1 _2016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3703_ _1250_ _1282_ _1281_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__o21ai_1
X_7471_ net395 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_1
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4683_ _2021_ _2083_ _2096_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__a21o_1
XFILLER_239_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6422_ _3128_ dmmu1.page_table\[0\]\[1\] _3135_ _3139_ vssd1 vssd1 vccd1 vccd1 _0536_
+ sky130_fd_sc_hd__a31o_1
X_3634_ _0917_ _1216_ _0920_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__a21o_1
XFILLER_146_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6353_ _3097_ vssd1 vssd1 vccd1 vccd1 _3098_ sky130_fd_sc_hd__buf_2
X_3565_ dmmu1.page_table\[8\]\[9\] dmmu1.page_table\[9\]\[9\] _0856_ vssd1 vssd1 vccd1
+ vccd1 _1149_ sky130_fd_sc_hd__mux2_1
XFILLER_115_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5425__A net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5304_ _1926_ _2479_ vssd1 vssd1 vccd1 vccd1 _2481_ sky130_fd_sc_hd__nor2_1
XFILLER_142_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6284_ _3053_ dmmu1.page_table\[5\]\[12\] _3037_ _3055_ vssd1 vssd1 vccd1 vccd1 _0482_
+ sky130_fd_sc_hd__a31o_1
X_3496_ _1080_ _1081_ _0881_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5235_ _2437_ _2438_ _1911_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__o21a_1
XFILLER_276_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6610__CLK clknet_leaf_53_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4150__C1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5166_ _2384_ dmmu0.page_table\[9\]\[2\] _2392_ vssd1 vssd1 vccd1 vccd1 _2395_ sky130_fd_sc_hd__and3_1
XFILLER_271_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4117_ immu_1.page_table\[0\]\[5\] immu_1.page_table\[1\]\[5\] _1448_ vssd1 vssd1
+ vccd1 vccd1 _1626_ sky130_fd_sc_hd__mux2_1
XFILLER_244_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5097_ _1922_ _2351_ vssd1 vssd1 vccd1 vccd1 _2352_ sky130_fd_sc_hd__or2_1
XANTENNA__5160__A _2216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6442__A1 _1898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4048_ _1456_ _1554_ _1558_ _1441_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__o211a_1
XANTENNA__6760__CLK clknet_leaf_0_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ _2793_ _2881_ vssd1 vssd1 vccd1 vccd1 _2885_ sky130_fd_sc_hd__and2_1
XANTENNA__7116__CLK clknet_leaf_30_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3819__S net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3559__A2 _1128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3716__C1 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5335__A _1933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input168_A c1_o_req_addr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input335_A ic1_mem_data[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input29_A c0_o_mem_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_46_core_clock clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_200_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4414__A _1373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5944__S _2848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5245__A _2370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3350_ _0869_ _0939_ _0941_ _0855_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__o211a_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ net123 vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__inv_6
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7460__A net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _1935_ _2302_ vssd1 vssd1 vccd1 vccd1 _2305_ sky130_fd_sc_hd__and2_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4295__S _1407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6076__A _2931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_85_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_281_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6424__A1 _3128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4308__B _1812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6971_ clknet_leaf_90_core_clock _0232_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[11\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7139__CLK clknet_leaf_33_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3212__B _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5922_ _2834_ dmmu0.page_table\[5\]\[5\] _2832_ vssd1 vssd1 vccd1 vccd1 _2839_ sky130_fd_sc_hd__and3_1
XFILLER_281_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4450__A3 _1924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5853_ net204 vssd1 vssd1 vccd1 vccd1 _2797_ sky130_fd_sc_hd__buf_2
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4804_ _2000_ _2170_ vssd1 vssd1 vccd1 vccd1 _2171_ sky130_fd_sc_hd__nor2_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4199__C1 _1360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5784_ _2749_ dmmu0.page_table\[13\]\[3\] _2751_ vssd1 vssd1 vccd1 vccd1 _2755_ sky130_fd_sc_hd__and3_1
XFILLER_221_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7289__CLK clknet_leaf_93_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4735_ _2014_ _2120_ _2129_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__a21o_1
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7454_ net58 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_1
XFILLER_135_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4666_ _1996_ _2083_ _2087_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__a21o_1
X_6405_ _1910_ vssd1 vssd1 vccd1 vccd1 _3128_ sky130_fd_sc_hd__buf_4
X_3617_ net121 _1199_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__or2_1
XANTENNA__5163__A1 _2211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7385_ net353 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_1
X_4597_ _2038_ immu_1.page_table\[13\]\[9\] _2032_ vssd1 vssd1 vccd1 vccd1 _2043_
+ sky130_fd_sc_hd__and3_1
XANTENNA__4697__C _2103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5155__A _2384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6336_ _3085_ dmmu1.page_table\[3\]\[6\] _3077_ _3087_ vssd1 vssd1 vccd1 vccd1 _0502_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__4910__A1 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3548_ _1129_ _1130_ _1131_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__and3_1
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6267_ _3042_ dmmu1.page_table\[5\]\[4\] _3038_ _3046_ vssd1 vssd1 vccd1 vccd1 _0474_
+ sky130_fd_sc_hd__a31o_1
XFILLER_170_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3479_ net151 dmmu1.long_off_reg\[1\] vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__xor2_1
XFILLER_95_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5218_ _2251_ _2408_ _2424_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__a21o_1
XFILLER_88_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6198_ _2994_ dmmu1.page_table\[7\]\[2\] _3000_ _3005_ vssd1 vssd1 vccd1 vccd1 _0446_
+ sky130_fd_sc_hd__a31o_1
XFILLER_276_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5149_ _2247_ _2369_ _2383_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__a21o_1
XFILLER_229_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5721__B1_N net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4977__A1 _1987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6506__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6433__B _3137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4729__A1 _2008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6194__A3 _3000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5049__B _2322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input285_A ic0_mem_data[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3792__B _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5154__A1 _2251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5065__A _2300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4901__A1 _2230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4480__B_N net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3313__A _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6185__A3 _2980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output671_A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5393__A1 _2531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5674__S _2690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3983__A _1442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7455__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4520_ net198 vssd1 vssd1 vccd1 vccd1 _1989_ sky130_fd_sc_hd__buf_4
XANTENNA__5145__A1 _2243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4451_ net99 vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__buf_4
X_3402_ _0958_ _0991_ _0899_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__o21a_1
X_7170_ clknet_leaf_35_core_clock _0431_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4382_ _0813_ _1883_ _1884_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__nor3_4
X_6121_ _1993_ _2943_ vssd1 vssd1 vccd1 vccd1 _2958_ sky130_fd_sc_hd__and2_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3333_ net19 _0924_ _0925_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__or3_1
XFILLER_285_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6052_ _2914_ dmmu1.page_table\[11\]\[10\] _2901_ _2916_ vssd1 vssd1 vccd1 vccd1
+ _0389_ sky130_fd_sc_hd__a31o_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3264_ _0856_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__buf_6
XFILLER_100_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5003_ _2284_ immu_1.page_table\[15\]\[9\] _2282_ vssd1 vssd1 vccd1 vccd1 _2293_
+ sky130_fd_sc_hd__and3_1
XFILLER_239_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4319__A _1584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3554__S1 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3195_ mem_dcache_arb.select _0810_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__nor2_1
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3223__A _0832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6529__CLK clknet_leaf_41_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4959__A1 _1987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6954_ clknet_leaf_82_core_clock _0215_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_241_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5620__A2 _2650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5905_ _2819_ dmmu0.page_table\[6\]\[12\] _2813_ vssd1 vssd1 vccd1 vccd1 _2828_ sky130_fd_sc_hd__and3_1
XFILLER_201_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6885_ clknet_leaf_84_core_clock _0146_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6679__CLK clknet_leaf_56_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5836_ _1958_ vssd1 vssd1 vccd1 vccd1 _2784_ sky130_fd_sc_hd__clkbuf_4
XFILLER_210_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6176__A3 _2981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4989__A _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5767_ _2736_ dmmu0.page_table\[4\]\[10\] _2731_ vssd1 vssd1 vccd1 vccd1 _2744_ sky130_fd_sc_hd__and3_1
XANTENNA__3893__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7506_ net393 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_1
X_4718_ _1959_ _2117_ vssd1 vssd1 vccd1 vccd1 _2118_ sky130_fd_sc_hd__or2_4
XFILLER_212_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5698_ _2682_ dmmu0.page_table\[2\]\[2\] _2702_ vssd1 vssd1 vccd1 vccd1 _2705_ sky130_fd_sc_hd__and3_1
X_4649_ _2072_ immu_1.page_table\[11\]\[6\] _2068_ vssd1 vssd1 vccd1 vccd1 _2076_
+ sky130_fd_sc_hd__and3_1
XFILLER_190_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7437_ net66 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3698__A1 _1279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7368_ net292 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_2
XFILLER_122_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6319_ _3076_ vssd1 vssd1 vccd1 vccd1 _3077_ sky130_fd_sc_hd__clkbuf_4
XFILLER_277_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7299_ clknet_leaf_44_core_clock _0560_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[8\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5332__B _2388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3870__A1 _1391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input200_A c1_sr_bus_data_o[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5611__A2 _2650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6163__B _2983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input96_A c0_sr_bus_data_o[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4899__A _2229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5375__A1 _2517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5507__B _2593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3308__A net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput360 ic1_mem_data[7] vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_2
XFILLER_222_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput371 ic1_wb_adr[2] vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_1
XFILLER_236_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput382 ic1_wb_stb vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_1
Xinput393 inner_wb_i_dat[13] vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_6
XFILLER_208_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3978__A _1447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6354__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3951_ _0813_ _1412_ _1436_ _1464_ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__a31o_1
XFILLER_90_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6073__B _2924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6670_ clknet_leaf_2_core_clock _0740_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_188_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3882_ net253 _1399_ _1386_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__mux2_4
XFILLER_204_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5621_ _2655_ dmmu0.page_table\[15\]\[5\] _2652_ vssd1 vssd1 vccd1 vccd1 _2659_ sky130_fd_sc_hd__and3_1
XANTENNA__5366__A1 _2503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3917__S _1425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4602__A _2000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5552_ _2232_ _2623_ _2625_ immu_0.page_table\[1\]\[4\] vssd1 vssd1 vccd1 vccd1 _0180_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3472__S0 _0858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4503_ _1977_ _1970_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__and2_1
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5417__B _2543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5118__A1 _2363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5483_ _2576_ immu_0.page_table\[4\]\[8\] _2574_ _2585_ vssd1 vssd1 vccd1 vccd1 _0151_
+ sky130_fd_sc_hd__a31o_1
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3218__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5136__C _2373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4434_ _1923_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__buf_4
X_7222_ clknet_leaf_16_core_clock _0483_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7153_ clknet_leaf_30_core_clock _0414_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[9\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_259_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4365_ immu_1.page_table\[0\]\[10\] immu_1.page_table\[1\]\[10\] _1439_ vssd1 vssd1
+ vccd1 vccd1 _1869_ sky130_fd_sc_hd__mux2_1
XANTENNA__3652__S _0896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6104_ _2948_ dmmu1.page_table\[9\]\[3\] _2942_ _2949_ vssd1 vssd1 vccd1 vccd1 _0408_
+ sky130_fd_sc_hd__a31o_1
XFILLER_258_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3316_ _0908_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__buf_4
XFILLER_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7084_ clknet_leaf_93_core_clock _0345_ vssd1 vssd1 vccd1 vccd1 dmmu0.long_off_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4296_ _1419_ _1800_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__or2_1
XANTENNA__6248__B _3020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6035_ _2898_ dmmu1.page_table\[11\]\[2\] _2902_ _2907_ vssd1 vssd1 vccd1 vccd1 _0381_
+ sky130_fd_sc_hd__a31o_1
X_3247_ _0846_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_1
XFILLER_239_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3301__B1 _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6264__A _2795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6937_ clknet_leaf_82_core_clock _0198_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6868_ clknet_leaf_73_core_clock _0129_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[6\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5357__A1 _2503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5819_ _2762_ dmmu0.page_table\[3\]\[5\] _2769_ vssd1 vssd1 vccd1 vccd1 _2775_ sky130_fd_sc_hd__and3_1
XFILLER_210_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6799_ clknet_leaf_8_core_clock _0060_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[7\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5608__A _2443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4512__A _1983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5109__A1 _2347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4317__C1 _1516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6439__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5343__A _2300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input150_A c1_o_mem_high_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input248_A dcache_wb_adr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6844__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input11_A c0_o_instr_long_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6388__A3 _3116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6994__CLK clknet_leaf_4_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4406__B _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5060__A3 _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3737__S _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4020__A1 _1516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5952__S _2848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6312__A3 _3057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5520__A1 _2603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6349__A _2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output634_A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4150_ _1442_ _1655_ _1657_ _1456_ vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__o211a_1
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4081_ immu_1.page_table\[6\]\[4\] immu_1.page_table\[7\]\[4\] _1439_ vssd1 vssd1
+ vccd1 vccd1 _1591_ sky130_fd_sc_hd__mux2_1
XFILLER_95_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6481__C1 _1911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput190 c1_sr_bus_addr[3] vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_4
XFILLER_270_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4983_ _2281_ vssd1 vssd1 vccd1 vccd1 _2282_ sky130_fd_sc_hd__buf_2
XFILLER_224_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3220__B _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6722_ clknet_leaf_67_core_clock _0792_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3934_ net366 vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__buf_4
XFILLER_189_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinterconnect_inner_718 vssd1 vssd1 vccd1 vccd1 interconnect_inner_718/HI c0_i_core_int_sreg[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinterconnect_inner_729 vssd1 vssd1 vccd1 vccd1 interconnect_inner_729/HI c1_i_core_int_sreg[6]
+ sky130_fd_sc_hd__conb_1
X_3865_ net318 net372 _1360_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__mux2_2
X_6653_ clknet_leaf_39_core_clock _0723_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_5604_ _2640_ dmmu0.page_table\[12\]\[12\] _2633_ vssd1 vssd1 vccd1 vccd1 _2648_
+ sky130_fd_sc_hd__and3_1
XFILLER_164_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6584_ clknet_leaf_47_core_clock _0654_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3796_ _1349_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_43_core_clock_A clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6717__CLK clknet_leaf_63_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4562__A2 _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5535_ _2603_ immu_0.page_table\[2\]\[7\] _2607_ _2616_ vssd1 vssd1 vccd1 vccd1 _0172_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__3770__A0 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5466_ _2561_ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput620 net620 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[6] sky130_fd_sc_hd__buf_2
XFILLER_117_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput631 net631 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[15] sky130_fd_sc_hd__buf_2
XANTENNA__6303__A3 _3058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput642 net642 vssd1 vssd1 vccd1 vccd1 ic1_mem_ppl_submit sky130_fd_sc_hd__buf_2
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7205_ clknet_leaf_28_core_clock _0466_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[6\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_4417_ _1908_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput653 net653 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[15] sky130_fd_sc_hd__buf_2
Xoutput664 net664 vssd1 vssd1 vccd1 vccd1 inner_wb_8_burst sky130_fd_sc_hd__buf_2
XANTENNA__6259__A _2931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5397_ _2531_ immu_0.page_table\[7\]\[6\] _2525_ _2534_ vssd1 vssd1 vccd1 vccd1 _0116_
+ sky130_fd_sc_hd__a31o_1
Xoutput675 net675 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[19] sky130_fd_sc_hd__buf_2
XANTENNA__6867__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput686 net686 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[7] sky130_fd_sc_hd__buf_2
Xoutput697 net697 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[1] sky130_fd_sc_hd__buf_2
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4348_ _1430_ _1849_ _1851_ _1416_ vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__o211a_1
X_7136_ clknet_leaf_13_core_clock _0397_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input3_A c0_o_c_instr_page vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_274_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7067_ clknet_leaf_5_core_clock _0328_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[6\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4078__A1 _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4279_ _1782_ _1783_ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__or2b_1
X_6018_ _2895_ _2880_ vssd1 vssd1 vccd1 vccd1 _2896_ sky130_fd_sc_hd__and2_1
XFILLER_46_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3411__A _0855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3589__B1 _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6441__B _3136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input198_A c1_sr_bus_data_o[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5057__B _2322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input365_A ic1_wb_adr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input59_A c0_o_req_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3420__A_N net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5502__A1 _2588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4388__S _1390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6169__A _2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5073__A _1930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5801__A _2762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5569__A1 _2235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7172__CLK clknet_leaf_37_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5248__A _2447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3650_ _0901_ _1231_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__or2_1
XFILLER_158_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3427__S0 _0897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3581_ _1163_ _1164_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__nand2_1
XFILLER_173_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5682__S _2690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7463__A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3752__A0 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5320_ _1944_ _2482_ vssd1 vssd1 vccd1 vccd1 _2490_ sky130_fd_sc_hd__and2_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5251_ _2230_ _2442_ _2450_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__a21o_1
XANTENNA__6079__A _2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4202_ _1648_ _1649_ _1650_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__o21ai_2
X_5182_ _2247_ _2390_ _2403_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__a21o_1
XFILLER_244_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4133_ _1535_ _1636_ _1638_ _1640_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__a31o_1
XFILLER_3_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3930__S _1443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5711__A _2709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4064_ immu_0.page_table\[12\]\[4\] immu_0.page_table\[13\]\[4\] immu_0.page_table\[14\]\[4\]
+ immu_0.page_table\[15\]\[4\] _1409_ _1420_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__mux4_1
XFILLER_216_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4327__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3231__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4966_ _2275_ vssd1 vssd1 vccd1 vccd1 _2276_ sky130_fd_sc_hd__clkinv_2
XFILLER_269_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6705_ clknet_leaf_62_core_clock _0775_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3917_ immu_0.page_table\[10\]\[0\] immu_0.page_table\[11\]\[0\] _1425_ vssd1 vssd1
+ vccd1 vccd1 _1431_ sky130_fd_sc_hd__mux2_1
XFILLER_149_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4783__A2 _2155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4897_ _2227_ _2219_ _2228_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__a21o_1
XANTENNA__5158__A _2217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6636_ clknet_leaf_40_core_clock _0706_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3848_ _1377_ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__clkbuf_1
XFILLER_192_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4997__A _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5732__A1 _1974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6567_ clknet_leaf_50_core_clock _0637_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3779_ _1340_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4091__S0 _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3743__A0 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5518_ _2606_ vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__clkbuf_4
XFILLER_218_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6498_ _3180_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5449_ net100 _2559_ vssd1 vssd1 vccd1 vccd1 _2566_ sky130_fd_sc_hd__and2_1
Xoutput450 net450 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[29] sky130_fd_sc_hd__buf_2
Xoutput461 net461 vssd1 vssd1 vccd1 vccd1 c0_i_req_data_valid sky130_fd_sc_hd__buf_2
Xoutput472 net472 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[12] sky130_fd_sc_hd__buf_2
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput483 net483 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[8] sky130_fd_sc_hd__buf_2
XFILLER_120_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput494 net494 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[17] sky130_fd_sc_hd__buf_2
XANTENNA__7045__CLK clknet_leaf_36_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7119_ clknet_leaf_28_core_clock _0380_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5621__A _2655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7195__CLK clknet_leaf_27_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4237__A _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input113_A c1_o_instr_long_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_core_clock clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4223__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3795__B _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3431__C1 _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6171__B _2983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3982__B1 _1441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3316__A _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3750__S _1322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_75_core_clock clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_238_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6562__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7458__A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4820_ _2166_ immu_1.page_table\[2\]\[6\] _2174_ vssd1 vssd1 vccd1 vccd1 _2181_ sky130_fd_sc_hd__and3_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6081__B _2924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5962__A1 _2805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4751_ _2139_ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__buf_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4765__A2 _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3702_ _1250_ _1281_ _1282_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__or3_1
X_4682_ _2089_ immu_1.page_table\[10\]\[8\] _2086_ vssd1 vssd1 vccd1 vccd1 _2096_
+ sky130_fd_sc_hd__and3_1
X_7470_ net394 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_1
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6421_ net201 _3137_ vssd1 vssd1 vccd1 vccd1 _3139_ sky130_fd_sc_hd__and2_1
X_3633_ dmmu0.page_table\[8\]\[10\] dmmu0.page_table\[9\]\[10\] dmmu0.page_table\[10\]\[10\]
+ dmmu0.page_table\[11\]\[10\] _0895_ net16 vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__mux4_1
XFILLER_174_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5714__A1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5706__A _2681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3564_ _0868_ _1147_ _0872_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__a21o_1
X_6352_ _2784_ _2170_ vssd1 vssd1 vccd1 vccd1 _3097_ sky130_fd_sc_hd__nor2_1
XANTENNA__4610__A _2038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_255_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7068__CLK clknet_leaf_4_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5425__B _2543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5303_ _2479_ vssd1 vssd1 vccd1 vccd1 _2480_ sky130_fd_sc_hd__clkbuf_4
X_6283_ net200 _3039_ vssd1 vssd1 vccd1 vccd1 _3055_ sky130_fd_sc_hd__and2_1
X_3495_ dmmu1.page_table\[0\]\[7\] dmmu1.page_table\[1\]\[7\] dmmu1.page_table\[2\]\[7\]
+ dmmu1.page_table\[3\]\[7\] _0858_ _0861_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__mux4_1
XFILLER_142_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3226__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5144__C _2373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5234_ net96 _2433_ _2427_ _2434_ net201 vssd1 vssd1 vccd1 vccd1 _2438_ sky130_fd_sc_hd__a32o_1
XFILLER_124_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5165_ _2224_ _2390_ _2394_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__a21o_1
XANTENNA__5493__A3 _2591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5441__A _1897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4116_ _1456_ _1620_ _1622_ _1624_ _1553_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__o221a_1
XFILLER_84_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5096_ _2295_ _2350_ vssd1 vssd1 vccd1 vccd1 _2351_ sky130_fd_sc_hd__or2_4
XFILLER_110_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5160__B _2388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4047_ _1555_ _1556_ _1557_ _1447_ _1451_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__a221o_1
XFILLER_209_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4453__A1 _1911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3896__A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6272__A _2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _2561_ vssd1 vssd1 vccd1 vccd1 _2884_ sky130_fd_sc_hd__buf_4
XFILLER_169_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4949_ _1977_ _2257_ _2265_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__a21o_1
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5705__A1 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6619_ clknet_leaf_53_core_clock _0689_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4064__S0 _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4520__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5335__B _2497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6130__A1 _2223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3570__S _1146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input230_A dcache_wb_4_burst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6585__CLK clknet_leaf_46_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input328_A ic0_wb_stb vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4444__A1 _1911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6182__A _2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5944__A1 _1933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4414__B net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5526__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4430__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output547_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _0869_ _0870_ _0872_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__o21a_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6928__CLK clknet_leaf_58_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5475__A3 _2574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5899__C _2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4683__A1 _2021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6970_ clknet_leaf_90_core_clock _0231_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5921_ _2232_ _2830_ _2838_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__a21o_1
XFILLER_253_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5852_ _2618_ dmmu1.page_table\[15\]\[3\] _2787_ _2796_ vssd1 vssd1 vccd1 vccd1 _0309_
+ sky130_fd_sc_hd__a31o_1
X_4803_ net190 net189 _1959_ vssd1 vssd1 vccd1 vccd1 _2170_ sky130_fd_sc_hd__or3_4
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5783_ _2226_ _2748_ _2754_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__a21o_1
XFILLER_221_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4734_ _2121_ immu_1.page_table\[6\]\[5\] _2123_ vssd1 vssd1 vccd1 vccd1 _2129_ sky130_fd_sc_hd__and3_1
XFILLER_159_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7453_ net75 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_1
XFILLER_119_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4665_ _2072_ immu_1.page_table\[10\]\[0\] _2086_ vssd1 vssd1 vccd1 vccd1 _2087_
+ sky130_fd_sc_hd__and3_1
XFILLER_147_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5436__A _1925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6404_ _3112_ dmmu1.page_table\[1\]\[8\] _3116_ _3127_ vssd1 vssd1 vccd1 vccd1 _0530_
+ sky130_fd_sc_hd__a31o_1
X_3616_ dmmu1.page_table\[12\]\[10\] dmmu1.page_table\[13\]\[10\] net120 vssd1 vssd1
+ vccd1 vccd1 _1199_ sky130_fd_sc_hd__mux2_1
XANTENNA__5163__A2 _2390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7384_ net342 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_2
XANTENNA__6360__A1 _3101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4596_ _2021_ _2030_ _2042_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__a21o_1
XFILLER_134_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6335_ net206 _3079_ vssd1 vssd1 vccd1 vccd1 _3087_ sky130_fd_sc_hd__and2_1
XFILLER_162_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3547_ _1129_ _1130_ _1131_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4910__A2 _2219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6112__A1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6266_ _2797_ _3040_ vssd1 vssd1 vccd1 vccd1 _3046_ sky130_fd_sc_hd__and2_1
X_3478_ _0880_ _1064_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__nand2_2
XFILLER_249_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5217_ _2416_ dmmu0.page_table\[8\]\[11\] _2410_ vssd1 vssd1 vccd1 vccd1 _2424_ sky130_fd_sc_hd__and3_1
X_6197_ _2793_ _3002_ vssd1 vssd1 vccd1 vccd1 _3005_ sky130_fd_sc_hd__and2_1
XFILLER_257_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5148_ _2371_ dmmu0.page_table\[10\]\[9\] _2373_ vssd1 vssd1 vccd1 vccd1 _2383_ sky130_fd_sc_hd__and3_1
XFILLER_56_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5079_ _2332_ immu_0.page_table\[12\]\[3\] _2336_ _2341_ vssd1 vssd1 vccd1 vccd1
+ _0800_ sky130_fd_sc_hd__a31o_1
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4977__A2 _2274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4515__A _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7233__CLK clknet_leaf_26_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4729__A2 _2120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3565__S _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5346__A _1944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4888__C _2221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input180_A c1_o_req_ppl_submit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4250__A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input278_A ic0_mem_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4901__A2 _2219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input41_A c0_o_mem_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6177__A _2891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5917__A1 _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output497_A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6600__CLK clknet_leaf_56_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output664_A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5256__A _2447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6342__A1 _3085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5145__A2 _2369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4450_ _1911_ immu_0.page_table\[11\]\[3\] _1924_ _1936_ vssd1 vssd1 vccd1 vccd1
+ _0576_ sky130_fd_sc_hd__a31o_1
XFILLER_171_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_48_core_clock_A clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_116_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3401_ _0989_ _0990_ _0906_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__mux2_1
X_4381_ _1874_ _1878_ _1882_ _1440_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__a31o_1
XANTENNA__7471__A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6120_ _2948_ dmmu1.page_table\[9\]\[11\] _2941_ _2957_ vssd1 vssd1 vccd1 vccd1 _0416_
+ sky130_fd_sc_hd__a31o_1
X_3332_ net46 net45 net48 net47 vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__or4_1
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5448__A3 _2557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4105__B1 _1613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6051_ _2895_ _2903_ vssd1 vssd1 vccd1 vccd1 _2916_ sky130_fd_sc_hd__and2_1
XANTENNA__6087__A _1991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3263_ net120 vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__buf_4
XFILLER_58_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7106__CLK clknet_leaf_32_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4656__A1 _2023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3504__A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5002_ _1985_ _2280_ _2292_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__a21o_1
XFILLER_39_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3194_ _0815_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_1
XFILLER_78_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4959__A2 _2257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6953_ clknet_leaf_84_core_clock _0214_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_121_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5081__A1 _2332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5904_ net94 _2811_ _2827_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__a21o_1
XFILLER_179_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6884_ clknet_leaf_84_core_clock _0145_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5835_ net95 _2766_ _2783_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__a21o_1
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3919__B1 _1432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5766_ _1948_ _2730_ _2743_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__a21o_1
XFILLER_194_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7505_ net392 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3395__A1 dmmu0.page_table\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4717_ net190 net189 vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__or2b_1
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5697_ _2224_ _2700_ _2704_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__a21o_1
XANTENNA__5166__A _2384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7436_ net59 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_1
XFILLER_135_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4648_ _2014_ _2066_ _2075_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__a21o_1
XFILLER_107_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7367_ net291 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_2
XFILLER_162_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4579_ _1996_ _2030_ _2033_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__a21o_1
XFILLER_146_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7381__A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6318_ _3075_ vssd1 vssd1 vccd1 vccd1 _3076_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_249_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7298_ clknet_leaf_43_core_clock _0559_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6249_ _3026_ dmmu1.page_table\[6\]\[11\] _3018_ _3034_ vssd1 vssd1 vccd1 vccd1 _0468_
+ sky130_fd_sc_hd__a31o_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_50_core_clock_A clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5072__A1 _2332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6623__CLK clknet_leaf_54_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6460__A _2971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input395_A inner_wb_i_dat[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3386__A1 _0963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input89_A c0_sr_bus_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5076__A _1933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4335__B1 _1432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7129__CLK clknet_leaf_29_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput350 ic1_mem_data[27] vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_2
Xinput361 ic1_mem_data[8] vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_2
XFILLER_48_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3310__A1 dmmu0.page_table\[1\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput372 ic1_wb_adr[3] vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_1
XFILLER_282_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput383 ic1_wb_we vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_1
Xinput394 inner_wb_i_dat[14] vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_6
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3978__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6354__B _3098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4155__A _1457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3950_ _1439_ _1441_ _1458_ _1463_ _0812_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__o221a_1
XFILLER_204_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3881_ net323 net377 _1390_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__mux2_1
XFILLER_231_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7466__A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5620_ _2233_ _2650_ _2658_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__a21o_1
XFILLER_176_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5366__A2 immu_0.page_table\[8\]\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5551_ _2229_ _2623_ _2625_ immu_0.page_table\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 _0179_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__4602__B _2045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3472__S1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4502_ net204 vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__buf_6
X_5482_ net103 _2577_ vssd1 vssd1 vccd1 vccd1 _2585_ sky130_fd_sc_hd__and2_1
X_7221_ clknet_leaf_27_core_clock _0482_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[5\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3218__B _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4433_ _1914_ _1922_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__or2_1
XFILLER_132_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7152_ clknet_leaf_33_core_clock _0413_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[9\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4364_ _1496_ _1867_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__or2_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6103_ _2795_ _2944_ vssd1 vssd1 vccd1 vccd1 _2949_ sky130_fd_sc_hd__and2_1
X_3315_ net16 vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__inv_2
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4295_ immu_0.page_table\[12\]\[9\] immu_0.page_table\[13\]\[9\] _1407_ vssd1 vssd1
+ vccd1 vccd1 _1800_ sky130_fd_sc_hd__mux2_1
X_7083_ clknet_leaf_5_core_clock _0344_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[5\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3234__A _0838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3246_ net128 net23 _0840_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__mux2_2
XFILLER_140_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6034_ _2793_ _2904_ vssd1 vssd1 vccd1 vccd1 _2907_ sky130_fd_sc_hd__and2_1
XFILLER_100_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3301__A1 _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6646__CLK clknet_leaf_42_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4991__C _2282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6264__B _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5054__A1 _2316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6936_ clknet_leaf_77_core_clock _0197_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6796__CLK clknet_leaf_10_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6867_ clknet_leaf_71_core_clock _0128_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_222_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6280__A _2931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5818_ _2232_ _2767_ _2774_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__a21o_1
XFILLER_179_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6798_ clknet_leaf_10_core_clock _0059_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[7\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3368__A1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5608__B _2296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4512__B _1970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5749_ _2223_ _2730_ _2734_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__a21o_1
XFILLER_182_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3409__A _0872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7419_ net389 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_1
XFILLER_163_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6439__B _3136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input143_A c1_o_mem_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5293__A1 _2245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input310_A ic0_wb_adr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5045__A1 _2316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4406__C net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4703__A _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3359__A1 dmmu0.page_table\[3\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3319__A _0901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6519__CLK clknet_leaf_36_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5534__A net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4323__A3 _1818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6349__B _2170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output627_A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4080_ _1496_ _1589_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__or2_1
XFILLER_283_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5284__A1 _2233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_255_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3295__B1 _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput180 c1_o_req_ppl_submit vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput191 c1_sr_bus_addr[4] vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5700__C _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4982_ _2084_ _2278_ vssd1 vssd1 vccd1 vccd1 _2281_ sky130_fd_sc_hd__or2_1
XFILLER_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6721_ clknet_leaf_63_core_clock _0791_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_251_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3933_ _1446_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5709__A _2709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinterconnect_inner_719 vssd1 vssd1 vccd1 vccd1 interconnect_inner_719/HI c0_i_core_int_sreg[10]
+ sky130_fd_sc_hd__conb_1
X_6652_ clknet_leaf_38_core_clock _0722_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3864_ _1387_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_1
X_5603_ _2251_ _2631_ _2647_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__a21o_1
XFILLER_137_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6000__A3 _2878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6583_ clknet_leaf_42_core_clock _0653_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3795_ net226 _1348_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__and2_1
XANTENNA__3229__A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5534_ net102 _2609_ vssd1 vssd1 vccd1 vccd1 _2616_ sky130_fd_sc_hd__and2_1
XFILLER_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5465_ _2562_ immu_0.page_table\[4\]\[0\] _2574_ _2575_ vssd1 vssd1 vccd1 vccd1 _0143_
+ sky130_fd_sc_hd__a31o_1
Xoutput610 net610 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[11] sky130_fd_sc_hd__buf_2
XFILLER_172_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput621 net621 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[7] sky130_fd_sc_hd__buf_2
XFILLER_145_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7204_ clknet_leaf_23_core_clock _0465_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[6\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput632 net632 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[1] sky130_fd_sc_hd__buf_2
X_4416_ _1373_ net388 vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__and2_1
Xoutput643 net643 vssd1 vssd1 vccd1 vccd1 ic1_mem_req sky130_fd_sc_hd__buf_2
Xoutput654 net654 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[1] sky130_fd_sc_hd__buf_2
Xoutput665 net665 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[0] sky130_fd_sc_hd__buf_2
X_5396_ _1942_ _2527_ vssd1 vssd1 vccd1 vccd1 _2534_ sky130_fd_sc_hd__and2_1
Xoutput676 net676 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[1] sky130_fd_sc_hd__buf_2
Xoutput687 net687 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[8] sky130_fd_sc_hd__buf_2
X_7135_ clknet_leaf_34_core_clock _0396_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput698 net698 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[2] sky130_fd_sc_hd__buf_2
X_4347_ _1423_ _1850_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__or2_1
XFILLER_113_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7066_ clknet_leaf_10_core_clock _0327_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[6\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4278_ net10 immu_0.high_addr_off\[5\] vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__or2_1
XFILLER_274_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4078__A2 _1582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3899__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6017_ net198 vssd1 vssd1 vccd1 vccd1 _2895_ sky130_fd_sc_hd__buf_2
X_3229_ net219 _0835_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__and2_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5610__C _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5027__A1 _2301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_core_clock clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3589__A1 _0901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6919_ clknet_leaf_75_core_clock _0180_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5619__A _2655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4523__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5354__A _1929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4896__C _2221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6811__CLK clknet_leaf_85_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input260_A dcache_wb_o_dat[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input358_A ic1_mem_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6169__B _2983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5073__B _2334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6230__A3 _3019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3748__S _1322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4433__A _1914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3427__S1 _0902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3580_ net154 dmmu1.long_off_reg\[4\] vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__or2_1
XFILLER_127_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5264__A _2447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5250_ _2447_ dmmu0.page_table\[7\]\[3\] _2445_ vssd1 vssd1 vccd1 vccd1 _2450_ sky130_fd_sc_hd__and3_1
XFILLER_114_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6297__A3 _3058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6079__B _2924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4201_ net8 immu_0.high_addr_off\[3\] vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__or2_1
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5181_ _2400_ dmmu0.page_table\[9\]\[9\] _2392_ vssd1 vssd1 vccd1 vccd1 _2403_ sky130_fd_sc_hd__and3_1
XFILLER_268_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4132_ _1479_ _1639_ _1434_ vssd1 vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__a21o_1
XFILLER_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5257__A1 _2240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4608__A _2038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4063_ immu_0.page_table\[8\]\[4\] immu_0.page_table\[9\]\[4\] immu_0.page_table\[10\]\[4\]
+ immu_0.page_table\[11\]\[4\] _1409_ _1420_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__mux4_1
XFILLER_283_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3231__B _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4965_ _2190_ _2273_ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__nand2_1
XFILLER_251_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3658__S _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5439__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6704_ clknet_leaf_45_core_clock _0774_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[15\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3916_ _1419_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__buf_4
X_4896_ _2204_ dmmu0.page_table\[0\]\[2\] _2221_ vssd1 vssd1 vccd1 vccd1 _2228_ sky130_fd_sc_hd__and3_1
XFILLER_177_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5158__B _2388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6635_ clknet_leaf_40_core_clock _0705_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3991__A1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3847_ _1373_ net259 vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__and2_4
XFILLER_285_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6834__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6566_ clknet_leaf_49_core_clock _0636_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3778_ net536 _1338_ _1339_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__and3b_2
XANTENNA__4091__S1 _1570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5517_ _1929_ _2605_ vssd1 vssd1 vccd1 vccd1 _2606_ sky130_fd_sc_hd__or2_1
XFILLER_285_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6497_ dmmu1.long_off_reg\[7\] _1983_ _3172_ vssd1 vssd1 vccd1 vccd1 _3180_ sky130_fd_sc_hd__mux2_1
XANTENNA__3393__S _0855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5174__A _2384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5448_ _2562_ immu_0.page_table\[5\]\[4\] _2557_ _2565_ vssd1 vssd1 vccd1 vccd1 _0136_
+ sky130_fd_sc_hd__a31o_1
Xoutput440 net440 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[1] sky130_fd_sc_hd__buf_2
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput451 net451 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[2] sky130_fd_sc_hd__buf_2
XANTENNA__5496__A1 _2588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput462 net462 vssd1 vssd1 vccd1 vccd1 c0_rst sky130_fd_sc_hd__buf_2
XANTENNA__6984__CLK clknet_leaf_7_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput473 net473 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[13] sky130_fd_sc_hd__buf_2
Xoutput484 net484 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[9] sky130_fd_sc_hd__buf_2
X_5379_ _2517_ immu_0.page_table\[8\]\[10\] _2509_ _2523_ vssd1 vssd1 vccd1 vccd1
+ _0109_ sky130_fd_sc_hd__a31o_1
XFILLER_154_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput495 net495 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[18] sky130_fd_sc_hd__buf_2
X_7118_ clknet_leaf_14_core_clock _0379_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3259__A0 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7049_ clknet_leaf_32_core_clock _0310_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4518__A _1987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3354__S0 _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4208__C1 _1432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A c1_o_c_data_page vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5420__A1 _2546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3982__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input71_A c0_o_req_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3734__A1 _0872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5084__A _1942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5487__A1 _2576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3345__S0 _0891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5250__C _2445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6707__CLK clknet_leaf_62_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6857__CLK clknet_leaf_69_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4750_ _2084_ _2136_ vssd1 vssd1 vccd1 vccd1 _2139_ sky130_fd_sc_hd__or2_1
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3701_ _1223_ _1225_ _1251_ _1248_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__a211oi_1
XFILLER_186_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4681_ _2019_ _2083_ _2095_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__a21o_1
XFILLER_119_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7474__A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6420_ _3128_ dmmu1.page_table\[0\]\[0\] _3135_ _3138_ vssd1 vssd1 vccd1 vccd1 _0535_
+ sky130_fd_sc_hd__a31o_1
X_3632_ _0901_ _1212_ _1214_ _0905_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__o211a_1
XANTENNA__5714__A2 _2700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3725__A1 _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6351_ _3095_ vssd1 vssd1 vccd1 vccd1 _3096_ sky130_fd_sc_hd__clkbuf_4
XFILLER_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3563_ dmmu1.page_table\[12\]\[9\] dmmu1.page_table\[13\]\[9\] _1146_ vssd1 vssd1
+ vccd1 vccd1 _1147_ sky130_fd_sc_hd__mux2_1
XFILLER_161_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5302_ _1922_ _2367_ vssd1 vssd1 vccd1 vccd1 _2479_ sky130_fd_sc_hd__or2_1
XFILLER_115_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6282_ _3053_ dmmu1.page_table\[5\]\[11\] _3037_ _3054_ vssd1 vssd1 vccd1 vccd1 _0481_
+ sky130_fd_sc_hd__a31o_1
XFILLER_255_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3494_ dmmu1.page_table\[4\]\[7\] dmmu1.page_table\[5\]\[7\] dmmu1.page_table\[6\]\[7\]
+ dmmu1.page_table\[7\]\[7\] _0892_ _0861_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__mux4_1
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3226__B _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3489__A0 _1072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5233_ _2223_ _2428_ _2436_ vssd1 vssd1 vccd1 vccd1 _2437_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4150__A1 _1442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5164_ _2384_ dmmu0.page_table\[9\]\[1\] _2392_ vssd1 vssd1 vccd1 vccd1 _2394_ sky130_fd_sc_hd__and3_1
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4115_ _1584_ _1623_ _1456_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__o21ai_1
XFILLER_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5095_ net83 net76 vssd1 vssd1 vccd1 vccd1 _2350_ sky130_fd_sc_hd__or2b_2
XFILLER_96_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6442__A3 _3134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4046_ immu_1.page_table\[4\]\[3\] immu_1.page_table\[5\]\[3\] _1443_ vssd1 vssd1
+ vccd1 vccd1 _1557_ sky130_fd_sc_hd__mux2_1
XFILLER_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_55_core_clock_A clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_271_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3896__B net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6272__B _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _2867_ dmmu1.page_table\[12\]\[1\] _2878_ _2883_ vssd1 vssd1 vccd1 vccd1 _0367_
+ sky130_fd_sc_hd__a31o_1
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4948_ _2262_ immu_1.page_table\[7\]\[4\] _2259_ vssd1 vssd1 vccd1 vccd1 _2265_ sky130_fd_sc_hd__and3_1
XFILLER_200_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4879_ net90 _1915_ vssd1 vssd1 vccd1 vccd1 _2213_ sky130_fd_sc_hd__or2_1
XFILLER_220_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6618_ clknet_leaf_53_core_clock _0688_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4801__A _2166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5705__A2 _2700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4064__S1 _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3716__A1 _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6549_ clknet_leaf_48_core_clock _0619_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_118_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5469__A1 _2576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7162__CLK clknet_leaf_11_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6130__A2 _2960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input223_A dcache_mem_o_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3652__A0 dmmu0.page_table\[6\]\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6182__B _2982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5807__A _2443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4711__A _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3327__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output442_A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4132__A1 _1479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_1_1_0_core_clock_A clknet_0_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4683__A2 _2083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3891__A0 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6424__A3 _3135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5632__A1 _2249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5688__S _2690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7469__A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5920_ _2834_ dmmu0.page_table\[5\]\[4\] _2832_ vssd1 vssd1 vccd1 vccd1 _2838_ sky130_fd_sc_hd__and3_1
XANTENNA__6373__A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_core_clock clknet_2_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_80_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5851_ _2795_ _2789_ vssd1 vssd1 vccd1 vccd1 _2796_ sky130_fd_sc_hd__and2_1
XFILLER_221_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4802_ _2025_ _2154_ _2169_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__a21o_1
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4199__B2 _1462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5782_ _2749_ dmmu0.page_table\[13\]\[2\] _2751_ vssd1 vssd1 vccd1 vccd1 _2754_ sky130_fd_sc_hd__and3_1
XANTENNA__7035__CLK clknet_leaf_12_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4733_ _2012_ _2120_ _2128_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__a21o_1
XFILLER_147_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5717__A _2709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4621__A _2054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7452_ net4 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_1
XFILLER_147_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4664_ _2085_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__buf_2
XFILLER_119_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5699__A1 _2227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6403_ net208 _3118_ vssd1 vssd1 vccd1 vccd1 _3127_ sky130_fd_sc_hd__and2_1
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3615_ dmmu1.page_table\[8\]\[10\] dmmu1.page_table\[9\]\[10\] dmmu1.page_table\[10\]\[10\]
+ dmmu1.page_table\[11\]\[10\] net120 net121 vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__mux4_1
XFILLER_266_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7383_ net331 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__clkbuf_2
X_4595_ _2038_ immu_1.page_table\[13\]\[8\] _2032_ vssd1 vssd1 vccd1 vccd1 _2042_
+ sky130_fd_sc_hd__and3_1
XANTENNA__7185__CLK clknet_leaf_13_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3237__A _0841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6334_ _3085_ dmmu1.page_table\[3\]\[5\] _3077_ _3086_ vssd1 vssd1 vccd1 vccd1 _0501_
+ sky130_fd_sc_hd__a31o_1
X_3546_ _1106_ _1108_ _1105_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__o21bai_1
XFILLER_135_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6265_ _3042_ dmmu1.page_table\[5\]\[3\] _3038_ _3045_ vssd1 vssd1 vccd1 vccd1 _0473_
+ sky130_fd_sc_hd__a31o_1
X_3477_ _1060_ _1063_ _0887_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__mux2_1
XFILLER_170_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5216_ _2249_ _2408_ _2423_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__a21o_1
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6196_ _2994_ dmmu1.page_table\[7\]\[1\] _3000_ _3004_ vssd1 vssd1 vccd1 vccd1 _0445_
+ sky130_fd_sc_hd__a31o_1
XFILLER_269_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5871__A1 _2805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5147_ _2245_ _2369_ _2382_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__a21o_1
XFILLER_84_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3882__A0 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5078_ _1935_ _2338_ vssd1 vssd1 vccd1 vccd1 _2341_ sky130_fd_sc_hd__and2_1
XFILLER_217_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7379__A clknet_leaf_19_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6283__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4029_ _1419_ _1539_ vssd1 vssd1 vccd1 vccd1 _1540_ sky130_fd_sc_hd__or2_1
XFILLER_231_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4515__B _1970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5627__A _2655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5346__B _2497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input173_A c1_o_req_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6458__A _2971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input340_A ic1_mem_data[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6177__B _2983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input34_A c0_o_mem_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3873__A0 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6193__A _2879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3610__A _0838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7058__CLK clknet_leaf_80_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5917__A2 _2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5393__A3 _2525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3756__S _1322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4441__A _1929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3400_ dmmu0.page_table\[12\]\[3\] dmmu0.page_table\[13\]\[3\] dmmu0.page_table\[14\]\[3\]
+ dmmu0.page_table\[15\]\[3\] _0898_ _0948_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__mux4_1
XANTENNA__5550__B1 _2625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4380_ _1874_ _1878_ _1882_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__a21oi_1
XFILLER_171_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3331_ net50 net49 net52 net51 vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__or4_1
XFILLER_124_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4105__A1 _1411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6050_ _2914_ dmmu1.page_table\[11\]\[9\] _2902_ _2915_ vssd1 vssd1 vccd1 vccd1 _0388_
+ sky130_fd_sc_hd__a31o_1
X_3262_ _0854_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__buf_4
X_5001_ _2284_ immu_1.page_table\[15\]\[8\] _2282_ vssd1 vssd1 vccd1 vccd1 _2292_
+ sky130_fd_sc_hd__and3_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3193_ net664 _0813_ net388 vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__and3_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5605__A1 _2253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6952_ clknet_leaf_82_core_clock _0213_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3711__S0 _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5903_ _2819_ dmmu0.page_table\[6\]\[11\] _2813_ vssd1 vssd1 vccd1 vccd1 _2827_ sky130_fd_sc_hd__and3_1
X_6883_ clknet_leaf_84_core_clock _0144_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5834_ _2777_ dmmu0.page_table\[3\]\[12\] _2768_ vssd1 vssd1 vccd1 vccd1 _2783_ sky130_fd_sc_hd__and3_1
XFILLER_201_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3919__A1 _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5765_ _2736_ dmmu0.page_table\[4\]\[9\] _2732_ vssd1 vssd1 vccd1 vccd1 _2743_ sky130_fd_sc_hd__and3_1
XANTENNA__4989__C _2282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5447__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4716_ _2025_ _2100_ _2116_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__a21o_1
X_7504_ net391 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4592__A1 _2016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5696_ _2682_ dmmu0.page_table\[2\]\[1\] _2702_ vssd1 vssd1 vccd1 vccd1 _2704_ sky130_fd_sc_hd__and3_1
XANTENNA__6575__CLK clknet_leaf_46_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7435_ clknet_opt_1_0_core_clock vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__buf_2
XFILLER_135_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4647_ _2072_ immu_1.page_table\[11\]\[5\] _2068_ vssd1 vssd1 vccd1 vccd1 _2075_
+ sky130_fd_sc_hd__and3_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7366_ net290 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_2
X_4578_ _2017_ immu_1.page_table\[13\]\[0\] _2032_ vssd1 vssd1 vccd1 vccd1 _2033_
+ sky130_fd_sc_hd__and3_1
XFILLER_150_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6317_ _2919_ _2193_ vssd1 vssd1 vccd1 vccd1 _3075_ sky130_fd_sc_hd__or2_1
X_3529_ dmmu1.page_table\[4\]\[8\] dmmu1.page_table\[5\]\[8\] dmmu1.page_table\[6\]\[8\]
+ dmmu1.page_table\[7\]\[8\] _0891_ _0860_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__mux4_1
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6278__A _2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7297_ clknet_leaf_43_core_clock _0558_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6097__A1 _2932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6248_ _1991_ _3020_ vssd1 vssd1 vccd1 vccd1 _3034_ sky130_fd_sc_hd__and2_1
XFILLER_249_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6179_ _2893_ _2983_ vssd1 vssd1 vccd1 vccd1 _2993_ sky130_fd_sc_hd__and2_1
XANTENNA__3855__A0 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7200__CLK clknet_leaf_22_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4526__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6021__A1 _2884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6918__CLK clknet_leaf_75_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5375__A3 _2510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4583__A1 _2008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3386__A2 _0967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input290_A ic0_mem_data[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4261__A _1523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input388_A inner_wb_err vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5076__B _2338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4335__A1 _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6188__A _2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6088__A1 _2932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5835__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput340 ic1_mem_data[18] vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__buf_2
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput351 ic1_mem_data[28] vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__buf_2
XFILLER_248_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput362 ic1_mem_data[9] vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_2
XFILLER_248_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput373 ic1_wb_adr[4] vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3941__S0 _1453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput384 inner_disable vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_4
Xinput395 inner_wb_i_dat[15] vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_6
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4436__A _1925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_4_0_core_clock_A clknet_2_2_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_251_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_opt_1_0_core_clock clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_opt_1_0_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_204_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3880_ _1398_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_1
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6598__CLK clknet_leaf_56_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5366__A3 _2510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5267__A _2458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5550_ _2226_ _2623_ _2625_ immu_0.page_table\[1\]\[2\] vssd1 vssd1 vccd1 vccd1 _0178_
+ sky130_fd_sc_hd__o22a_1
XFILLER_129_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4501_ _1898_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__buf_6
XFILLER_157_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5481_ _2576_ immu_0.page_table\[4\]\[7\] _2574_ _2584_ vssd1 vssd1 vccd1 vccd1 _0150_
+ sky130_fd_sc_hd__a31o_1
XFILLER_117_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5118__A3 _2353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7220_ clknet_leaf_27_core_clock _0481_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[5\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_117_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4432_ _1921_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__buf_6
XANTENNA__4326__B2 _1830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7151_ clknet_leaf_33_core_clock _0412_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6098__A _2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4363_ immu_1.page_table\[4\]\[10\] immu_1.page_table\[5\]\[10\] _1524_ vssd1 vssd1
+ vccd1 vccd1 _1867_ sky130_fd_sc_hd__mux2_1
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6102_ _2931_ vssd1 vssd1 vccd1 vccd1 _2948_ sky130_fd_sc_hd__buf_4
X_3314_ _0903_ _0904_ _0906_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__mux2_1
X_7082_ clknet_leaf_5_core_clock _0343_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[5\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_263_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4294_ immu_0.page_table\[14\]\[9\] immu_0.page_table\[15\]\[9\] _1408_ vssd1 vssd1
+ vccd1 vccd1 _1799_ sky130_fd_sc_hd__mux2_1
XFILLER_140_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6033_ _2898_ dmmu1.page_table\[11\]\[1\] _2902_ _2906_ vssd1 vssd1 vccd1 vccd1 _0380_
+ sky130_fd_sc_hd__a31o_1
X_3245_ _0845_ vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_core_clock clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3250__A _0848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6251__A1 _3026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6935_ clknet_leaf_58_core_clock _0196_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6866_ clknet_leaf_71_core_clock _0127_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5817_ _2762_ dmmu0.page_table\[3\]\[4\] _2769_ vssd1 vssd1 vccd1 vccd1 _2774_ sky130_fd_sc_hd__and3_1
XANTENNA__5357__A3 _2510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6797_ clknet_leaf_10_core_clock _0058_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5177__A _2400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4565__A1 _2021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3368__A2 _0944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5748_ _2709_ dmmu0.page_table\[4\]\[1\] _2732_ vssd1 vssd1 vccd1 vccd1 _2734_ sky130_fd_sc_hd__and3_1
XFILLER_210_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5109__A3 _2353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5679_ _2693_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7392__A net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5905__A _2819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4317__A1 _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7418_ net710 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_1
XFILLER_135_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7349_ net303 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_2
XFILLER_116_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_core_clock clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_249_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5640__A _1914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5293__A2 _2462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input136_A c1_o_mem_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input303_A ic0_mem_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_260_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6740__CLK clknet_leaf_66_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4005__A0 immu_1.page_table\[0\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6890__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5815__A _2762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7246__CLK clknet_leaf_26_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3335__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5520__A3 _2607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output522_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3819__A0 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5284__A2 _2462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput170 c1_o_req_addr[15] vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
XANTENNA__6365__B _3098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3295__A1 _0855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput181 c1_sr_bus_addr[0] vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_4
Xinput192 c1_sr_bus_addr[5] vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_1
XFILLER_236_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4166__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _2279_ vssd1 vssd1 vccd1 vccd1 _2280_ sky130_fd_sc_hd__clkbuf_4
XFILLER_224_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3932_ net367 vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__inv_2
XFILLER_211_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6720_ clknet_leaf_63_core_clock _0790_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4795__A1 _2019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6651_ clknet_leaf_38_core_clock _0721_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3863_ net247 _1385_ _1386_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__mux2_4
XFILLER_176_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5602_ _2640_ dmmu0.page_table\[12\]\[11\] _2633_ vssd1 vssd1 vccd1 vccd1 _2647_
+ sky130_fd_sc_hd__and3_1
X_6582_ clknet_leaf_45_core_clock _0652_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3794_ _0839_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__clkbuf_2
XFILLER_176_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5533_ _2603_ immu_0.page_table\[2\]\[6\] _2607_ _2615_ vssd1 vssd1 vccd1 vccd1 _0171_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__3229__B _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5464_ _1925_ _2573_ vssd1 vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__nor2_1
Xoutput600 net600 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[8] sky130_fd_sc_hd__buf_2
XFILLER_160_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput611 net611 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[12] sky130_fd_sc_hd__buf_2
XFILLER_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7203_ clknet_leaf_22_core_clock _0464_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput622 net622 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[8] sky130_fd_sc_hd__buf_2
X_4415_ _1907_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkbuf_1
Xoutput633 net633 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[2] sky130_fd_sc_hd__buf_2
X_5395_ _2531_ immu_0.page_table\[7\]\[5\] _2525_ _2533_ vssd1 vssd1 vccd1 vccd1 _0115_
+ sky130_fd_sc_hd__a31o_1
Xoutput644 net644 vssd1 vssd1 vccd1 vccd1 ic1_rst sky130_fd_sc_hd__buf_2
XANTENNA__6613__CLK clknet_leaf_54_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3245__A _0845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput655 net655 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[2] sky130_fd_sc_hd__buf_2
Xoutput666 net666 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[10] sky130_fd_sc_hd__buf_2
Xoutput677 net677 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[20] sky130_fd_sc_hd__buf_2
X_7134_ clknet_leaf_13_core_clock _0395_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput688 net688 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[9] sky130_fd_sc_hd__buf_2
X_4346_ immu_0.page_table\[2\]\[10\] immu_0.page_table\[3\]\[10\] _1407_ vssd1 vssd1
+ vccd1 vccd1 _1850_ sky130_fd_sc_hd__mux2_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput699 net699 vssd1 vssd1 vccd1 vccd1 inner_wb_o_dat[3] sky130_fd_sc_hd__buf_2
XFILLER_98_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7065_ clknet_leaf_11_core_clock _0326_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4277_ net10 immu_0.high_addr_off\[5\] vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__and2_1
X_6016_ _2884_ dmmu1.page_table\[12\]\[9\] _2878_ _2894_ vssd1 vssd1 vccd1 vccd1 _0375_
+ sky130_fd_sc_hd__a31o_1
XFILLER_246_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3228_ _0818_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__buf_4
XFILLER_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6763__CLK clknet_leaf_86_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4076__A _1584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7119__CLK clknet_leaf_28_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7387__A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4804__A _2000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6918_ clknet_leaf_75_core_clock _0179_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6849_ clknet_leaf_73_core_clock _0110_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5635__A _2370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_62_core_clock_A clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5354__B _2407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5502__A3 _2591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4710__A1 _2019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input253_A dcache_wb_adr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6466__A _2971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5370__A _1942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6463__A1 _1972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5801__C _2750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_253_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6215__A1 _3010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4433__B _1922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5726__A0 immu_1.high_addr_off\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5248__C _2445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3764__S _1322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4200_ net8 immu_0.high_addr_off\[3\] vssd1 vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__nand2_1
X_5180_ _2245_ _2390_ _2402_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__a21o_1
XANTENNA__6786__CLK clknet_leaf_0_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4131_ immu_0.page_table\[12\]\[6\] immu_0.page_table\[13\]\[6\] immu_0.page_table\[14\]\[6\]
+ immu_0.page_table\[15\]\[6\] _1601_ _1430_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__mux4_1
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5257__A2 _2442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4062_ immu_0.page_table\[4\]\[4\] immu_0.page_table\[5\]\[4\] immu_0.page_table\[6\]\[4\]
+ immu_0.page_table\[7\]\[4\] _1409_ _1420_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__mux4_1
XFILLER_56_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5711__C _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6206__A1 _2994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4964_ _2273_ vssd1 vssd1 vccd1 vccd1 _2274_ sky130_fd_sc_hd__buf_4
XFILLER_212_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6703_ clknet_leaf_45_core_clock _0773_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[15\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5439__B _2559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3915_ _1424_ _1428_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__nand2_1
X_4895_ _2226_ vssd1 vssd1 vccd1 vccd1 _2227_ sky130_fd_sc_hd__clkbuf_4
X_3846_ _1376_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_1
X_6634_ clknet_leaf_40_core_clock _0704_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6565_ clknet_leaf_49_core_clock _0635_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3777_ _0838_ _1168_ _1211_ _1279_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__or4_1
XFILLER_138_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4997__C _2282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5455__A _2310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5516_ net85 net84 _2317_ vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__or3_4
XANTENNA__4940__A1 _1995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6496_ _3179_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__clkbuf_1
X_5447_ net99 _2559_ vssd1 vssd1 vccd1 vccd1 _2565_ sky130_fd_sc_hd__and2_1
XFILLER_160_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput430 net430 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[10] sky130_fd_sc_hd__buf_2
Xoutput441 net441 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[20] sky130_fd_sc_hd__buf_2
Xoutput452 net452 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[30] sky130_fd_sc_hd__buf_2
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput463 net463 vssd1 vssd1 vccd1 vccd1 c1_clk sky130_fd_sc_hd__clkbuf_1
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput474 net474 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[14] sky130_fd_sc_hd__buf_2
X_5378_ _2314_ _2512_ vssd1 vssd1 vccd1 vccd1 _2523_ sky130_fd_sc_hd__and2_1
Xoutput485 net485 vssd1 vssd1 vccd1 vccd1 c1_i_mem_exception sky130_fd_sc_hd__buf_2
Xoutput496 net496 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[19] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_6_core_clock clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_core_clock
+ sky130_fd_sc_hd__clkbuf_16
X_7117_ clknet_leaf_30_core_clock _0378_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[12\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_259_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4329_ _1783_ _1785_ _1782_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__a21o_1
XFILLER_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5190__A _2217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5621__C _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7048_ clknet_leaf_37_core_clock _0309_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4518__B _1970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3354__S1 _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6509__CLK clknet_leaf_59_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4759__A1 _2010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4534__A _1999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7091__CLK clknet_leaf_2_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3982__A2 _1494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5184__A1 _2249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5365__A _1937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input370_A ic1_wb_adr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5084__B _2338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input64_A c0_o_req_addr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4709__A _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6436__A1 _1898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4998__A1 _1981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3345__S1 _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5962__A3 _2859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ net52 dmmu0.long_off_reg\[7\] vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4680_ _2089_ immu_1.page_table\[10\]\[7\] _2086_ vssd1 vssd1 vccd1 vccd1 _2095_
+ sky130_fd_sc_hd__and3_1
XANTENNA__5175__A1 _2240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3631_ _0908_ _1213_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__or2_1
XFILLER_186_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5275__A _2458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6350_ _3094_ vssd1 vssd1 vccd1 vccd1 _3095_ sky130_fd_sc_hd__dlymetal6s2s_1
X_3562_ _0856_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__buf_4
XFILLER_127_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4610__C _2049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5301_ _2253_ _2461_ _2478_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__a21o_1
XFILLER_255_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6281_ net199 _3039_ vssd1 vssd1 vccd1 vccd1 _3054_ sky130_fd_sc_hd__and2_1
XFILLER_142_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3493_ _1065_ _1069_ _1079_ _0819_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__o2bb2a_4
XFILLER_115_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7490__A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5232_ net201 _2430_ net408 vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__a21bo_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3489__A1 _1075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5163_ _2211_ _2390_ _2393_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__a21o_1
XANTENNA__4619__A _2054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4114_ immu_1.page_table\[14\]\[5\] immu_1.page_table\[15\]\[5\] _1438_ vssd1 vssd1
+ vccd1 vccd1 _1623_ sky130_fd_sc_hd__mux2_1
XFILLER_110_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5094_ _2347_ immu_0.page_table\[12\]\[10\] _2335_ _2349_ vssd1 vssd1 vccd1 vccd1
+ _0807_ sky130_fd_sc_hd__a31o_1
XFILLER_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4045_ _1448_ immu_1.page_table\[6\]\[3\] net367 vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__o21a_1
XFILLER_271_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4453__A3 _1924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _2791_ _2881_ vssd1 vssd1 vccd1 vccd1 _2883_ sky130_fd_sc_hd__and2_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4947_ _1974_ _2257_ _2264_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__a21o_1
XFILLER_177_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4878_ net83 net76 net85 net84 vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__or4_4
XFILLER_228_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6617_ clknet_leaf_62_core_clock _0687_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3829_ _1367_ vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_1
XFILLER_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5185__A _2400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6548_ clknet_leaf_48_core_clock _0618_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[13\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_229_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6479_ _1989_ _3156_ _3170_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__a21o_1
XFILLER_106_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7307__CLK clknet_leaf_19_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5913__A _2681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4529__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4444__A3 _1924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input216_A dcache_mem_o_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5807__B _2589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5823__A _2681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4439__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output435_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6409__A1 _3128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3891__A1 _1405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6824__CLK clknet_leaf_59_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6373__B _3098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4840__B1 _2192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5850_ net203 vssd1 vssd1 vccd1 vccd1 _2795_ sky130_fd_sc_hd__buf_2
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4801_ _2166_ immu_1.page_table\[4\]\[10\] _2156_ vssd1 vssd1 vccd1 vccd1 _2169_
+ sky130_fd_sc_hd__and3_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6974__CLK clknet_leaf_0_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5781_ _2223_ _2748_ _2753_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__a21o_1
XFILLER_221_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4902__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4732_ _2121_ immu_1.page_table\[6\]\[4\] _2123_ vssd1 vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__and3_1
XFILLER_147_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4663_ _2084_ _2081_ vssd1 vssd1 vccd1 vccd1 _2085_ sky130_fd_sc_hd__or2_1
X_7451_ net65 vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_1
XFILLER_174_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3518__A _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3614_ _1195_ _1196_ net122 vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__mux2_1
X_6402_ _3112_ dmmu1.page_table\[1\]\[7\] _3116_ _3126_ vssd1 vssd1 vccd1 vccd1 _0529_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__5699__A2 _2700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4594_ _2019_ _2030_ _2041_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__a21o_1
X_7382_ net408 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__clkbuf_1
XANTENNA__6360__A3 _3096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6333_ net205 _3079_ vssd1 vssd1 vccd1 vccd1 _3086_ sky130_fd_sc_hd__and2_1
X_3545_ net48 dmmu0.long_off_reg\[3\] vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__or2_1
XANTENNA__3952__S _0811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6264_ _2795_ _3040_ vssd1 vssd1 vccd1 vccd1 _3045_ sky130_fd_sc_hd__and2_1
XFILLER_170_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3476_ _1061_ _1062_ _0881_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__mux2_1
XANTENNA__6112__A3 _2942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5215_ _2416_ dmmu0.page_table\[8\]\[10\] _2410_ vssd1 vssd1 vccd1 vccd1 _2423_ sky130_fd_sc_hd__and3_1
XFILLER_142_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6195_ _2791_ _3002_ vssd1 vssd1 vccd1 vccd1 _3004_ sky130_fd_sc_hd__and2_1
XFILLER_229_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5146_ _2371_ dmmu0.page_table\[10\]\[8\] _2373_ vssd1 vssd1 vccd1 vccd1 _2382_ sky130_fd_sc_hd__and3_1
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3882__A1 _1399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5077_ _2332_ immu_0.page_table\[12\]\[2\] _2336_ _2340_ vssd1 vssd1 vccd1 vccd1
+ _0799_ sky130_fd_sc_hd__a31o_1
XFILLER_244_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4028_ immu_0.page_table\[12\]\[3\] immu_0.page_table\[13\]\[3\] _1407_ vssd1 vssd1
+ vccd1 vccd1 _1539_ sky130_fd_sc_hd__mux2_1
XFILLER_56_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3634__A1 _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5979_ _2867_ dmmu1.page_table\[13\]\[8\] _2859_ _2871_ vssd1 vssd1 vccd1 vccd1 _0361_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__7395__A net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3398__B1 _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4812__A _2166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5139__A1 _2233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input166_A c1_o_req_addr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6847__CLK clknet_leaf_69_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input333_A ic1_mem_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3873__A1 _1393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input27_A c0_o_mem_addr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6474__A _2190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6997__CLK clknet_leaf_62_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6193__B _3002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4722__A _2084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3484__S0 _0900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5256__C _2445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6342__A3 _3077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5550__A1 _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3772__S _0839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3330_ _0899_ _0907_ _0916_ _0922_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__o22a_1
XFILLER_112_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3261_ net122 vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__buf_4
XFILLER_98_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4169__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5000_ _1983_ _2280_ _2291_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__a21o_1
XFILLER_285_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3192_ _0814_ vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_1
XFILLER_285_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6384__A _3115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3801__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7002__CLK clknet_leaf_37_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6951_ clknet_leaf_84_core_clock _0212_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1_1_core_clock clknet_1_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_1_1_1_core_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5081__A3 _2336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5902_ _1950_ _2811_ _2826_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__a21o_1
XFILLER_281_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6882_ clknet_leaf_71_core_clock _0143_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3711__S1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5369__A1 _2517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5833_ net94 _2766_ _2782_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__a21o_1
XANTENNA__7152__CLK clknet_leaf_33_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4632__A _2000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5764_ _1946_ _2730_ _2742_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__a21o_1
XANTENNA__3475__S0 _0858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7503_ net390 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5447__B _2559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4715_ _2106_ immu_1.page_table\[9\]\[10\] _2102_ vssd1 vssd1 vccd1 vccd1 _2116_
+ sky130_fd_sc_hd__and3_1
XANTENNA__4592__A2 _2030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3395__A3 dmmu0.page_table\[3\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5695_ _2211_ _2700_ _2703_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__a21o_1
XANTENNA__3248__A _0839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5166__C _2392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7434_ net395 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_1
X_4646_ _2012_ _2066_ _2074_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__a21o_1
XFILLER_107_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4577_ _2031_ vssd1 vssd1 vccd1 vccd1 _2032_ sky130_fd_sc_hd__buf_2
X_7365_ net289 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_2
XFILLER_162_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3682__S _1146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6316_ _3069_ dmmu1.page_table\[4\]\[12\] _3057_ _3074_ vssd1 vssd1 vccd1 vccd1 _0495_
+ sky130_fd_sc_hd__a31o_1
XFILLER_1_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3528_ dmmu1.page_table\[0\]\[8\] dmmu1.page_table\[1\]\[8\] dmmu1.page_table\[2\]\[8\]
+ dmmu1.page_table\[3\]\[8\] _0891_ _0860_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__mux4_1
XFILLER_1_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7296_ clknet_leaf_44_core_clock _0557_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_226_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_core_clock clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_67_core_clock_A clknet_3_2_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_115_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6247_ _3026_ dmmu1.page_table\[6\]\[10\] _3018_ _3033_ vssd1 vssd1 vccd1 vccd1 _0467_
+ sky130_fd_sc_hd__a31o_1
X_3459_ _0913_ _1046_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__or2_1
XFILLER_103_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6178_ _2977_ dmmu1.page_table\[8\]\[8\] _2981_ _2992_ vssd1 vssd1 vccd1 vccd1 _0439_
+ sky130_fd_sc_hd__a31o_1
XFILLER_130_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5129_ _2372_ vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__clkbuf_4
XFILLER_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6294__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3430__B net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5072__A3 _2336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5638__A _1914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4542__A _1910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6460__C _3159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4583__A2 _2030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_84_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input283_A ic0_mem_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3592__S _1169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6188__B _2255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4099__A1 _1479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput330 ic1_mem_ack vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_1
XFILLER_282_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput341 ic1_mem_data[19] vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_2
Xinput352 ic1_mem_data[29] vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_2
XFILLER_208_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput363 ic1_wb_adr[0] vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4717__A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput374 ic1_wb_adr[5] vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3310__A3 dmmu0.page_table\[3\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput385 inner_embed_mode vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_6
XFILLER_152_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3941__S1 _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput396 inner_wb_i_dat[1] vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_16
XFILLER_208_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5599__A1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7175__CLK clknet_leaf_11_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4452__A _1937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4500_ _1939_ dmmu1.page_table\[14\]\[3\] _1964_ _1975_ vssd1 vssd1 vccd1 vccd1 _0587_
+ sky130_fd_sc_hd__a31o_1
X_5480_ net102 _2577_ vssd1 vssd1 vccd1 vccd1 _2584_ sky130_fd_sc_hd__and2_1
XFILLER_157_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4431_ _1917_ _1920_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__or2_2
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5523__A1 _2603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4326__A2 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6379__A _1910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5283__A _2458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3534__B1 _0854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7150_ clknet_leaf_35_core_clock _0411_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4362_ _1523_ _1865_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__or2_1
XFILLER_263_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6098__B _2944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6101_ _2932_ dmmu1.page_table\[9\]\[2\] _2942_ _2947_ vssd1 vssd1 vccd1 vccd1 _0407_
+ sky130_fd_sc_hd__a31o_1
X_3313_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__buf_4
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7081_ clknet_leaf_9_core_clock _0342_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[5\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4293_ _1424_ _1797_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__or2_1
XFILLER_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6032_ _2791_ _2904_ vssd1 vssd1 vccd1 vccd1 _2906_ sky130_fd_sc_hd__and2_1
X_3244_ net127 net22 _0840_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__mux2_1
XFILLER_246_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4627__A _2054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5054__A3 _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6934_ clknet_leaf_75_core_clock _0195_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6542__CLK clknet_leaf_48_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6865_ clknet_leaf_70_core_clock _0126_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4362__A _1523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5816_ _2229_ _2767_ _2773_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__a21o_1
X_6796_ clknet_leaf_10_core_clock _0057_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4565__A2 _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5747_ _2210_ _2730_ _2733_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__a21o_1
XANTENNA__5762__A1 _2242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6692__CLK clknet_leaf_42_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5678_ _2226_ immu_0.high_addr_off\[2\] _2690_ vssd1 vssd1 vccd1 vccd1 _2693_ sky130_fd_sc_hd__mux2_1
XFILLER_175_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7417_ clknet_leaf_92_core_clock vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__buf_2
XANTENNA__6289__A _3059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4629_ net189 net190 vssd1 vssd1 vccd1 vccd1 _2062_ sky130_fd_sc_hd__or2b_1
XFILLER_135_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3525__B1 _0957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7348_ net302 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_2
XANTENNA__7048__CLK clknet_leaf_37_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7279_ clknet_leaf_21_core_clock _0540_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_277_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5640__B _2215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4537__A _1961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input129_A c1_o_mem_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5045__A3 _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5368__A _1940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3439__S0 _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4703__C _2103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input94_A c0_sr_bus_data_o[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3764__A0 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5815__B dmmu0.page_table\[3\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6199__A _2795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3335__B net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3819__A1 _1361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6481__A2 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput160 c1_o_mem_sel[0] vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__buf_2
XFILLER_248_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput171 c1_o_req_addr[1] vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_2
Xinput182 c1_sr_bus_addr[10] vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6565__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput193 c1_sr_bus_addr[6] vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_1
XFILLER_263_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4980_ _1999_ _2278_ vssd1 vssd1 vccd1 vccd1 _2279_ sky130_fd_sc_hd__nor2_1
XFILLER_251_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3931_ _1442_ _1444_ vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__and2_1
XANTENNA__4795__A2 _2155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6650_ clknet_leaf_39_core_clock _0720_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5709__C _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3862_ _0811_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__buf_6
XFILLER_258_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5601_ _2249_ _2631_ _2646_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__a21o_1
XFILLER_149_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6581_ clknet_leaf_46_core_clock _0651_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[10\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3793_ _1347_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_1
XANTENNA__7493__A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5532_ net101 _2609_ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__and2_1
XFILLER_157_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5463_ _2573_ vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__clkbuf_4
XFILLER_172_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput601 net601 vssd1 vssd1 vccd1 vccd1 ic0_mem_addr[9] sky130_fd_sc_hd__buf_2
XFILLER_105_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7202_ clknet_leaf_15_core_clock _0463_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput612 net612 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[13] sky130_fd_sc_hd__buf_2
X_4414_ _1373_ net387 vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__and2_1
Xoutput623 net623 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[9] sky130_fd_sc_hd__buf_2
Xoutput634 net634 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[3] sky130_fd_sc_hd__buf_2
X_5394_ _1940_ _2527_ vssd1 vssd1 vccd1 vccd1 _2533_ sky130_fd_sc_hd__and2_1
XFILLER_132_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput645 net645 vssd1 vssd1 vccd1 vccd1 ic1_wb_ack sky130_fd_sc_hd__buf_2
Xoutput656 net656 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[3] sky130_fd_sc_hd__buf_2
Xoutput667 net667 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[11] sky130_fd_sc_hd__buf_2
XANTENNA__4180__B1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7133_ clknet_leaf_14_core_clock _0394_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput678 net678 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[21] sky130_fd_sc_hd__buf_2
X_4345_ immu_0.page_table\[0\]\[10\] immu_0.page_table\[1\]\[10\] _1425_ vssd1 vssd1
+ vccd1 vccd1 _1849_ sky130_fd_sc_hd__mux2_1
XFILLER_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput689 net689 vssd1 vssd1 vccd1 vccd1 inner_wb_cyc sky130_fd_sc_hd__buf_2
XFILLER_259_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7064_ clknet_leaf_10_core_clock _0325_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4276_ _1755_ _1781_ _1569_ net243 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6908__CLK clknet_leaf_75_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6015_ _2893_ _2881_ vssd1 vssd1 vccd1 vccd1 _2894_ sky130_fd_sc_hd__and2_1
X_3227_ _0834_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4357__A _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3261__A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5680__A0 _2229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5027__A3 _2298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4476__D_N net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6917_ clknet_leaf_58_core_clock _0178_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5983__A1 _2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3443__C1 _0855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4804__B _2170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4092__A _1408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5619__C _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6848_ clknet_leaf_69_core_clock _0109_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[8\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6779_ clknet_leaf_87_core_clock _0040_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3746__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5916__A _2834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4820__A _2166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3436__A _0863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4710__A2 _2101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3870__S _1386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6588__CLK clknet_leaf_45_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input246_A dcache_wb_adr[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5370__B _2512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6463__A2 _3157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4206__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3985__B1 _1497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5726__A1 _1995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5826__A _2777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4730__A _2121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6151__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5561__A _2190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4130_ _1478_ _1637_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__or2_1
XFILLER_268_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4061_ immu_0.page_table\[0\]\[4\] immu_0.page_table\[1\]\[4\] immu_0.page_table\[2\]\[4\]
+ immu_0.page_table\[3\]\[4\] _1409_ _1570_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__mux4_1
XFILLER_3_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4177__A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4608__C _2049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4963_ _1999_ _2272_ vssd1 vssd1 vccd1 vccd1 _2273_ sky130_fd_sc_hd__or2_1
X_6702_ clknet_leaf_45_core_clock _0772_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[15\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3914_ immu_0.page_table\[8\]\[0\] immu_0.page_table\[9\]\[0\] _1408_ vssd1 vssd1
+ vccd1 vccd1 _1428_ sky130_fd_sc_hd__mux2_1
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4894_ net97 vssd1 vssd1 vccd1 vccd1 _2226_ sky130_fd_sc_hd__buf_4
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6633_ clknet_leaf_40_core_clock _0703_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3845_ _1373_ net258 vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__and2_4
XANTENNA__3955__S _1425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3728__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4640__A _2054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6564_ clknet_leaf_49_core_clock _0634_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6390__A1 _3112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3776_ _1194_ _1228_ _1254_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__or3_1
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5455__B _2559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5226__B1_N net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5515_ _2603_ immu_0.page_table\[3\]\[10\] _2590_ _2604_ vssd1 vssd1 vccd1 vccd1
+ _0164_ sky130_fd_sc_hd__a31o_1
XFILLER_285_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4940__A2 _2257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6495_ dmmu1.long_off_reg\[6\] _1981_ _3172_ vssd1 vssd1 vccd1 vccd1 _3179_ sky130_fd_sc_hd__mux2_1
XANTENNA__3256__A _0851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5174__C _2392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5446_ _2562_ immu_0.page_table\[5\]\[3\] _2557_ _2564_ vssd1 vssd1 vccd1 vccd1 _0135_
+ sky130_fd_sc_hd__a31o_1
Xoutput420 net420 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[2] sky130_fd_sc_hd__buf_2
XANTENNA__6142__A1 _2242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput431 net431 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[11] sky130_fd_sc_hd__buf_2
XFILLER_160_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6730__CLK clknet_leaf_66_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput442 net442 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[21] sky130_fd_sc_hd__buf_2
XANTENNA__5496__A3 _2591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput453 net453 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[31] sky130_fd_sc_hd__buf_2
Xoutput464 net464 vssd1 vssd1 vccd1 vccd1 c1_disable sky130_fd_sc_hd__buf_2
XFILLER_259_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput475 net475 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[15] sky130_fd_sc_hd__buf_2
X_5377_ _2517_ immu_0.page_table\[8\]\[9\] _2510_ _2522_ vssd1 vssd1 vccd1 vccd1 _0108_
+ sky130_fd_sc_hd__a31o_1
XFILLER_160_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput486 net486 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[0] sky130_fd_sc_hd__buf_2
X_7116_ clknet_leaf_30_core_clock _0377_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[12\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput497 net497 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[1] sky130_fd_sc_hd__buf_2
XFILLER_113_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4328_ net11 immu_0.high_addr_off\[6\] vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__or2_1
XFILLER_101_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input1_A c0_o_c_data_page vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5190__B _2407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7047_ clknet_leaf_37_core_clock _0308_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_274_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4259_ _1523_ _1764_ _1530_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__o21ai_1
XFILLER_274_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6880__CLK clknet_leaf_70_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3664__C1 _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7398__A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_255_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4208__A1 _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4759__A2 _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5420__A3 _2541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5708__A1 _2240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3865__S _1360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5646__A _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4550__A _1977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6381__A1 _3112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input196_A c1_sr_bus_addr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4392__A0 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5365__B _2512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input363_A ic1_wb_adr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input57_A c0_o_mem_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4447__A1 _1911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4998__A2 _2280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3655__C1 _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6603__CLK clknet_leaf_41_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3958__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3630_ dmmu0.page_table\[14\]\[10\] dmmu0.page_table\[15\]\[10\] net15 vssd1 vssd1
+ vccd1 vccd1 _1213_ sky130_fd_sc_hd__mux2_1
XANTENNA__6372__A1 _3101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5175__A2 _2390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3561_ _0859_ _1144_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__and2_1
XFILLER_255_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5300_ _2473_ dmmu0.page_table\[14\]\[12\] _2463_ vssd1 vssd1 vccd1 vccd1 _2478_
+ sky130_fd_sc_hd__and3_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6280_ _2931_ vssd1 vssd1 vccd1 vccd1 _3053_ sky130_fd_sc_hd__clkbuf_4
X_3492_ _0929_ _1076_ _1078_ _0957_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__a22o_1
XFILLER_154_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5231_ _2432_ _2435_ _1911_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__o21a_1
XANTENNA__7109__CLK clknet_leaf_32_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6387__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5291__A _2370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5162_ _2384_ dmmu0.page_table\[9\]\[0\] _2392_ vssd1 vssd1 vccd1 vccd1 _2393_ sky130_fd_sc_hd__and3_1
XFILLER_271_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4113_ _1581_ _1621_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__nor2_1
XFILLER_96_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5093_ _2314_ _2338_ vssd1 vssd1 vccd1 vccd1 _2349_ sky130_fd_sc_hd__and2_1
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4438__A1 _1911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7259__CLK clknet_leaf_25_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4044_ immu_1.page_table\[7\]\[3\] _1448_ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__or2b_1
XFILLER_244_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5938__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5995_ _2867_ dmmu1.page_table\[12\]\[0\] _2878_ _2882_ vssd1 vssd1 vccd1 vccd1 _0366_
+ sky130_fd_sc_hd__a31o_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3949__B1 _1462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4946_ _2262_ immu_1.page_table\[7\]\[3\] _2259_ vssd1 vssd1 vccd1 vccd1 _2264_ sky130_fd_sc_hd__and3_1
XFILLER_220_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4877_ _2210_ vssd1 vssd1 vccd1 vccd1 _2211_ sky130_fd_sc_hd__buf_4
XFILLER_177_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5466__A _2561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4370__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6616_ clknet_leaf_54_core_clock _0686_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3828_ _1363_ net265 vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__and2_1
XFILLER_137_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5185__B dmmu0.page_table\[9\]\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6547_ clknet_leaf_51_core_clock _0617_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[13\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3759_ _1329_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6478_ _2190_ immu_1.page_table\[8\]\[10\] _3158_ vssd1 vssd1 vccd1 vccd1 _3170_
+ sky130_fd_sc_hd__and3_1
XFILLER_279_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5469__A3 _2574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4126__B1 _1614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5429_ _2312_ _2543_ vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__and2_1
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4677__A1 _2014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3714__A net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6626__CLK clknet_leaf_56_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4545__A _1910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input111_A c1_o_instr_long_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input209_A c1_sr_bus_data_o[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5929__A1 _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_74_core_clock_A clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6776__CLK clknet_leaf_85_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3595__S _1169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5376__A _2312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4711__C _2103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6106__A1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4668__A1 _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4455__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4840__A1 _1974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4800_ _2023_ _2155_ _2168_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__a21o_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5780_ _2749_ dmmu0.page_table\[13\]\[1\] _2751_ vssd1 vssd1 vccd1 vccd1 _2753_ sky130_fd_sc_hd__and3_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4731_ _2010_ _2120_ _2127_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__a21o_1
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7450_ net64 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__clkbuf_1
X_4662_ _1998_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__clkbuf_4
XFILLER_266_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4621__C _2049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6401_ net207 _3118_ vssd1 vssd1 vccd1 vccd1 _3126_ sky130_fd_sc_hd__and2_1
XFILLER_174_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3613_ dmmu1.page_table\[4\]\[10\] dmmu1.page_table\[5\]\[10\] dmmu1.page_table\[6\]\[10\]
+ dmmu1.page_table\[7\]\[10\] net120 net121 vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__mux4_1
X_7381_ net408 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_1
X_4593_ _2038_ immu_1.page_table\[13\]\[7\] _2032_ vssd1 vssd1 vccd1 vccd1 _2041_
+ sky130_fd_sc_hd__and3_1
XFILLER_134_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6332_ _2931_ vssd1 vssd1 vccd1 vccd1 _3085_ sky130_fd_sc_hd__buf_4
X_3544_ net48 dmmu0.long_off_reg\[3\] vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__nand2_1
XFILLER_155_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_35_core_clock clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6263_ _3042_ dmmu1.page_table\[5\]\[2\] _3038_ _3044_ vssd1 vssd1 vccd1 vccd1 _0472_
+ sky130_fd_sc_hd__a31o_1
X_3475_ dmmu1.page_table\[8\]\[6\] dmmu1.page_table\[9\]\[6\] dmmu1.page_table\[10\]\[6\]
+ dmmu1.page_table\[11\]\[6\] _0858_ _0861_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__mux4_1
XFILLER_115_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5214_ _2247_ _2409_ _2422_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__a21o_1
XANTENNA__7081__CLK clknet_leaf_9_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6194_ _2994_ dmmu1.page_table\[7\]\[0\] _3000_ _3003_ vssd1 vssd1 vccd1 vccd1 _0444_
+ sky130_fd_sc_hd__a31o_1
X_5145_ _2243_ _2369_ _2381_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__a21o_1
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _1933_ _2338_ vssd1 vssd1 vccd1 vccd1 _2340_ sky130_fd_sc_hd__and2_1
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4027_ immu_0.page_table\[14\]\[3\] immu_0.page_table\[15\]\[3\] _1408_ vssd1 vssd1
+ vccd1 vccd1 _1538_ sky130_fd_sc_hd__mux2_1
XFILLER_37_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _1985_ _2861_ vssd1 vssd1 vccd1 vccd1 _2871_ sky130_fd_sc_hd__and2_1
XFILLER_212_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3398__A1 _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4929_ _2237_ dmmu0.page_table\[0\]\[11\] _2220_ vssd1 vssd1 vccd1 vccd1 _2252_ sky130_fd_sc_hd__and3_1
XANTENNA__5196__A _2400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_core_clock clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6336__A1 _3085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5139__A2 _2369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5627__C _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5924__A _2834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6458__C _3159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input159_A c1_o_mem_req vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input326_A ic0_wb_sel[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5075__A1 _2332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4722__B _2118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3484__S1 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4214__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6327__A1 _3069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4889__A1 _2211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5834__A _2777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5550__A2 _2623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3260_ _0853_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_2
XFILLER_239_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3191_ net664 _0813_ net387 vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__and3_1
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6941__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3801__B _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6950_ clknet_leaf_81_core_clock _0211_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4813__A1 _2008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5901_ _2819_ dmmu0.page_table\[6\]\[10\] _2813_ vssd1 vssd1 vccd1 vccd1 _2826_ sky130_fd_sc_hd__and3_1
XFILLER_241_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6881_ clknet_leaf_71_core_clock _0142_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[5\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7496__A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5832_ _2777_ dmmu0.page_table\[3\]\[11\] _2768_ vssd1 vssd1 vccd1 vccd1 _2782_ sky130_fd_sc_hd__and3_1
XFILLER_222_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5369__A2 immu_0.page_table\[8\]\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4913__A _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5763_ _2736_ dmmu0.page_table\[4\]\[8\] _2732_ vssd1 vssd1 vccd1 vccd1 _2742_ sky130_fd_sc_hd__and3_1
XANTENNA__4632__B _2064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7502_ net404 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3475__S1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4714_ _2023_ _2101_ _2115_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__a21o_1
XFILLER_147_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5694_ _2682_ dmmu0.page_table\[2\]\[0\] _2702_ vssd1 vssd1 vccd1 vccd1 _2703_ sky130_fd_sc_hd__and3_1
XFILLER_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7433_ net394 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_1
X_4645_ _2072_ immu_1.page_table\[11\]\[4\] _2068_ vssd1 vssd1 vccd1 vccd1 _2074_
+ sky130_fd_sc_hd__and3_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5744__A _2443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7364_ net287 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_2
X_4576_ _1999_ _2028_ vssd1 vssd1 vccd1 vccd1 _2031_ sky130_fd_sc_hd__or2_1
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6315_ net200 _3059_ vssd1 vssd1 vccd1 vccd1 _3074_ sky130_fd_sc_hd__and2_1
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3527_ _1087_ _1088_ _1095_ _1112_ vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__a31o_4
X_7295_ clknet_leaf_44_core_clock _0556_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3264__A _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6246_ _2895_ _3020_ vssd1 vssd1 vccd1 vccd1 _3033_ sky130_fd_sc_hd__and2_1
XANTENNA__6097__A3 _2942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3458_ dmmu0.page_table\[8\]\[5\] dmmu0.page_table\[9\]\[5\] _0896_ vssd1 vssd1 vccd1
+ vccd1 _1046_ sky130_fd_sc_hd__mux2_1
XFILLER_103_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6177_ _2891_ _2983_ vssd1 vssd1 vccd1 vccd1 _2992_ sky130_fd_sc_hd__and2_1
Xclkbuf_2_2_0_core_clock clknet_1_1_1_core_clock vssd1 vssd1 vccd1 vccd1 clknet_2_2_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
X_3389_ _0977_ _0978_ _0855_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__mux2_1
X_5128_ _2216_ _2367_ vssd1 vssd1 vccd1 vccd1 _2372_ sky130_fd_sc_hd__or2_1
XFILLER_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6294__B _3060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5059_ _1944_ _2322_ vssd1 vssd1 vccd1 vccd1 _2329_ sky130_fd_sc_hd__and2_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4823__A _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6021__A3 _2877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5638__B _2217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3240__A0 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3873__S _1386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5654__A _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input276_A ic0_mem_ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput320 ic0_wb_adr[5] vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__buf_2
XANTENNA__3902__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput331 ic1_mem_data[0] vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput342 ic1_mem_data[1] vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_1
XFILLER_248_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput353 ic1_mem_data[2] vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_2
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput364 ic1_wb_adr[10] vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_2
XANTENNA__5048__A1 _2316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput375 ic1_wb_adr[6] vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput386 inner_ext_irq vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_1
XFILLER_275_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput397 inner_wb_i_dat[2] vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_8
XFILLER_263_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4209__S _1425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5599__A2 _2632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4452__B _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5220__A1 _2253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3349__A _0863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4430_ net710 _1919_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__or2_1
XFILLER_144_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3534__A1 _0869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4361_ immu_1.page_table\[6\]\[10\] immu_1.page_table\[7\]\[10\] _1524_ vssd1 vssd1
+ vccd1 vccd1 _1865_ sky130_fd_sc_hd__mux2_1
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6100_ _2793_ _2944_ vssd1 vssd1 vccd1 vccd1 _2947_ sky130_fd_sc_hd__and2_1
XFILLER_113_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3312_ net17 vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__buf_4
XFILLER_112_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7080_ clknet_leaf_11_core_clock _0341_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[5\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4292_ immu_0.page_table\[10\]\[9\] immu_0.page_table\[11\]\[9\] _1425_ vssd1 vssd1
+ vccd1 vccd1 _1797_ sky130_fd_sc_hd__mux2_1
X_6031_ _2898_ dmmu1.page_table\[11\]\[0\] _2902_ _2905_ vssd1 vssd1 vccd1 vccd1 _0379_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__6395__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3243_ _0844_ vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_1
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4908__A _2105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4119__S _1448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6251__A3 _3018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6933_ clknet_leaf_57_core_clock _0194_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_281_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4643__A _2072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6864_ clknet_leaf_71_core_clock _0125_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_222_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5815_ _2762_ dmmu0.page_table\[3\]\[3\] _2769_ vssd1 vssd1 vccd1 vccd1 _2773_ sky130_fd_sc_hd__and3_1
XFILLER_195_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6795_ clknet_leaf_80_core_clock _0056_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6837__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5177__C _2392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5746_ _2709_ dmmu0.page_table\[4\]\[0\] _2732_ vssd1 vssd1 vccd1 vccd1 _2733_ sky130_fd_sc_hd__and3_1
XANTENNA__5762__A2 _2730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4970__B1 _2277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5677_ _2692_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5474__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7416_ net211 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_1
X_4628_ _2025_ _2046_ _2061_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__a21o_1
XFILLER_135_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6987__CLK clknet_leaf_7_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7347_ net299 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_2
XFILLER_104_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4559_ _2016_ _2002_ _2018_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__a21o_1
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7278_ clknet_leaf_21_core_clock _0539_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5278__A1 _2224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6229_ _2793_ _3021_ vssd1 vssd1 vccd1 vccd1 _3024_ sky130_fd_sc_hd__and2_1
XFILLER_249_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4818__A _2166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4537__B _1998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4238__C1 _1535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_13_core_clock_A clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__5450__A1 _2562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4553__A _1979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5368__B _2512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3439__S1 _0864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input393_A inner_wb_i_dat[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input87_A c0_sr_bus_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5384__A _1930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6199__B _3002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7142__CLK clknet_leaf_29_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4728__A _2121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput150 c1_o_mem_high_addr[0] vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_2
XFILLER_283_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput161 c1_o_mem_sel[1] vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput172 c1_o_req_addr[2] vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput183 c1_sr_bus_addr[11] vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_1
Xinput194 c1_sr_bus_addr[7] vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7292__CLK clknet_leaf_43_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5559__A _1929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3930_ immu_1.page_table\[6\]\[0\] immu_1.page_table\[7\]\[0\] _1443_ vssd1 vssd1
+ vccd1 vccd1 _1444_ sky130_fd_sc_hd__mux2_1
XFILLER_189_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3861_ net317 net371 _1360_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__mux2_2
XFILLER_149_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5600_ _2640_ dmmu0.page_table\[12\]\[10\] _2633_ vssd1 vssd1 vccd1 vccd1 _2646_
+ sky130_fd_sc_hd__and3_1
XFILLER_258_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6580_ clknet_leaf_49_core_clock _0650_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[10\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3792_ net225 _0993_ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__and2_1
XFILLER_176_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5531_ _2603_ immu_0.page_table\[2\]\[5\] _2607_ _2614_ vssd1 vssd1 vccd1 vccd1 _0170_
+ sky130_fd_sc_hd__a31o_1
XFILLER_145_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5294__A _2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3807__A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5462_ _1929_ _2572_ vssd1 vssd1 vccd1 vccd1 _2573_ sky130_fd_sc_hd__or2_1
XFILLER_274_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7201_ clknet_leaf_15_core_clock _0462_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput602 net602 vssd1 vssd1 vccd1 vccd1 ic0_mem_cache_flush sky130_fd_sc_hd__buf_2
X_4413_ _1906_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__clkbuf_2
Xoutput613 net613 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[14] sky130_fd_sc_hd__buf_2
Xoutput624 net624 vssd1 vssd1 vccd1 vccd1 ic1_clk sky130_fd_sc_hd__clkbuf_1
X_5393_ _2531_ immu_0.page_table\[7\]\[4\] _2525_ _2532_ vssd1 vssd1 vccd1 vccd1 _0114_
+ sky130_fd_sc_hd__a31o_1
Xoutput635 net635 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[4] sky130_fd_sc_hd__buf_2
XFILLER_160_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_0_0_core_clock_A clknet_2_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput646 net646 vssd1 vssd1 vccd1 vccd1 ic1_wb_err sky130_fd_sc_hd__buf_2
X_7132_ clknet_leaf_34_core_clock _0393_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput657 net657 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[4] sky130_fd_sc_hd__buf_2
XFILLER_132_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput668 net668 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[12] sky130_fd_sc_hd__buf_2
XFILLER_259_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4344_ _1430_ _1847_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__or2_1
Xoutput679 net679 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[22] sky130_fd_sc_hd__buf_2
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7063_ clknet_leaf_10_core_clock _0324_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4638__A _2054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4275_ _1579_ _1761_ _1780_ inner_wb_arbiter.o_sel_sig vssd1 vssd1 vccd1 vccd1 _1781_
+ sky130_fd_sc_hd__a31o_1
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6014_ net209 vssd1 vssd1 vccd1 vccd1 _2893_ sky130_fd_sc_hd__buf_2
X_3226_ net218 _0824_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__and2_1
XFILLER_239_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_4_core_clock_A clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5432__A1 _2546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6916_ clknet_leaf_74_core_clock _0177_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3994__A1 _1424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6847_ clknet_leaf_69_core_clock _0108_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[8\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6778_ clknet_leaf_85_core_clock _0039_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_79_core_clock_A clknet_3_3_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_139_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7015__CLK clknet_leaf_11_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5729_ _2722_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7165__CLK clknet_leaf_10_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5932__A _2834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4548__A _1910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6466__C _3159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3357__S0 _0898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input141_A c1_o_mem_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input239_A dcache_wb_adr[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__A1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3737__A1 _1317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6003__A _2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output458_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5842__A _1995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6532__CLK clknet_leaf_46_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4458__A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4060_ _1430_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__buf_4
XFILLER_49_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6682__CLK clknet_leaf_41_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6206__A3 _3000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5289__A _2458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4962_ net188 net181 net190 net189 vssd1 vssd1 vccd1 vccd1 _2272_ sky130_fd_sc_hd__or4_4
XFILLER_269_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7038__CLK clknet_leaf_9_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6701_ clknet_leaf_42_core_clock _0771_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3913_ _1424_ _1426_ _1416_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__a21oi_1
X_4893_ _2224_ _2219_ _2225_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__a21o_1
X_6632_ clknet_leaf_41_core_clock _0702_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3844_ _1375_ vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_1
XFILLER_177_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3728__A1 _0854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6563_ clknet_leaf_49_core_clock _0633_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3775_ _1337_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_1
XFILLER_164_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5514_ net93 _2593_ vssd1 vssd1 vccd1 vccd1 _2604_ sky130_fd_sc_hd__and2_1
XFILLER_157_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6494_ _3178_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__clkbuf_1
X_5445_ net98 _2559_ vssd1 vssd1 vccd1 vccd1 _2564_ sky130_fd_sc_hd__and2_1
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput410 net410 vssd1 vssd1 vccd1 vccd1 c0_i_mc_core_int sky130_fd_sc_hd__buf_2
XANTENNA__6142__A2 _2960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput421 net421 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[3] sky130_fd_sc_hd__buf_2
XFILLER_218_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput432 net432 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[12] sky130_fd_sc_hd__buf_2
XANTENNA__5752__A _2681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput443 net443 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[22] sky130_fd_sc_hd__buf_2
XFILLER_172_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5376_ _2312_ _2512_ vssd1 vssd1 vccd1 vccd1 _2522_ sky130_fd_sc_hd__and2_1
Xoutput454 net454 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[3] sky130_fd_sc_hd__buf_2
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput465 net465 vssd1 vssd1 vccd1 vccd1 c1_i_core_int_sreg[0] sky130_fd_sc_hd__buf_2
Xoutput476 net476 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[1] sky130_fd_sc_hd__buf_2
X_7115_ clknet_leaf_30_core_clock _0376_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[12\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput487 net487 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[10] sky130_fd_sc_hd__buf_2
XANTENNA__3361__C1 _0918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput498 net498 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[20] sky130_fd_sc_hd__buf_2
X_4327_ net11 immu_0.high_addr_off\[6\] vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__nand2_1
XFILLER_160_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3272__A _0857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_259_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7046_ clknet_leaf_32_core_clock _0307_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4258_ immu_1.page_table\[10\]\[8\] immu_1.page_table\[11\]\[8\] _1493_ vssd1 vssd1
+ vccd1 vccd1 _1764_ sky130_fd_sc_hd__mux2_1
XFILLER_86_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5653__A1 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3209_ _0825_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_1
X_4189_ immu_1.page_table\[8\]\[7\] immu_1.page_table\[9\]\[7\] _1443_ vssd1 vssd1
+ vccd1 vccd1 _1696_ sky130_fd_sc_hd__mux2_1
XFILLER_227_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5405__A1 _2531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4208__A2 _1712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4307__S _1453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3511__S0 _0897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4831__A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5708__A2 _2700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_259_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4392__A1 _1892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input189_A c1_sr_bus_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6555__CLK clknet_leaf_50_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3881__S _1390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5662__A _2682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input356_A ic1_mem_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5892__A1 _2235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4278__A net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4709__C _2103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6436__A3 _3135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3910__A _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4217__S _1407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5837__A _2784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3186__A2 _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3560_ dmmu1.page_table\[14\]\[9\] dmmu1.page_table\[15\]\[9\] _0856_ vssd1 vssd1
+ vccd1 vccd1 _1144_ sky130_fd_sc_hd__mux2_1
XANTENNA__5275__C _2464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_core_clock clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_127_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3491_ _1055_ _1077_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5230_ net92 _2433_ _2427_ _2434_ net197 vssd1 vssd1 vccd1 vccd1 _2435_ sky130_fd_sc_hd__a32o_1
XFILLER_154_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6387__B _3118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5883__A1 _2223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5161_ _2391_ vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4619__C _2049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4112_ immu_1.page_table\[12\]\[5\] immu_1.page_table\[13\]\[5\] _1493_ vssd1 vssd1
+ vccd1 vccd1 _1621_ sky130_fd_sc_hd__mux2_1
XFILLER_110_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5092_ _2347_ immu_0.page_table\[12\]\[9\] _2336_ _2348_ vssd1 vssd1 vccd1 vccd1
+ _0806_ sky130_fd_sc_hd__a31o_1
XFILLER_229_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7499__A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4043_ immu_1.page_table\[0\]\[3\] immu_1.page_table\[1\]\[3\] immu_1.page_table\[2\]\[3\]
+ immu_1.page_table\[3\]\[3\] _1453_ _1454_ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__mux4_1
XFILLER_284_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4916__A _2242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3646__A0 _1211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3820__A _1362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4127__S _1601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5994_ _2879_ _2881_ vssd1 vssd1 vccd1 vccd1 _2882_ sky130_fd_sc_hd__and2_1
XFILLER_252_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3949__A1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4945_ _1972_ _2257_ _2263_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__a21o_1
XFILLER_220_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4651__A _2072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4876_ net92 vssd1 vssd1 vccd1 vccd1 _2210_ sky130_fd_sc_hd__buf_6
XFILLER_220_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6578__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3827_ _1366_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_1
XFILLER_220_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6615_ clknet_leaf_53_core_clock _0685_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3267__A _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6546_ clknet_leaf_50_core_clock _0616_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[13\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3758_ net149 net44 _1322_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__mux2_2
XFILLER_116_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6477_ _1987_ _3157_ _3169_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__a21o_1
X_3689_ dmmu1.page_table\[2\]\[11\] dmmu1.page_table\[3\]\[11\] _0856_ vssd1 vssd1
+ vccd1 vccd1 _1271_ sky130_fd_sc_hd__mux2_1
XANTENNA__5482__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5428_ _2546_ immu_0.page_table\[6\]\[8\] _2541_ _2552_ vssd1 vssd1 vccd1 vccd1 _0129_
+ sky130_fd_sc_hd__a31o_1
XFILLER_279_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4677__A2 _2083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5359_ _1928_ _2512_ vssd1 vssd1 vccd1 vccd1 _2513_ sky130_fd_sc_hd__and2_1
XANTENNA__3885__A0 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7203__CLK clknet_leaf_22_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5626__A1 _2243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7029_ clknet_leaf_7_core_clock _0290_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[13\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4037__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5929__A2 _2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input104_A c0_sr_bus_data_o[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3876__S _1386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4561__A _2017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5376__B _2512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5392__A _1937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3905__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4668__A2 _2083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3876__A0 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6409__A3 _3115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3971__S0 _1453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4736__A _2121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4840__A2 _2189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6720__CLK clknet_leaf_63_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4471__A _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4730_ _2121_ immu_1.page_table\[6\]\[3\] _2123_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__and3_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4661_ _2082_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__clkbuf_4
XFILLER_202_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6400_ _3112_ dmmu1.page_table\[1\]\[6\] _3116_ _3125_ vssd1 vssd1 vccd1 vccd1 _0528_
+ sky130_fd_sc_hd__a31o_1
XFILLER_174_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3612_ dmmu1.page_table\[0\]\[10\] dmmu1.page_table\[1\]\[10\] dmmu1.page_table\[2\]\[10\]
+ dmmu1.page_table\[3\]\[10\] net120 net121 vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__mux4_1
XFILLER_266_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5553__B1 _2625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7380_ net407 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_1
X_4592_ _2016_ _2030_ _2040_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__a21o_1
XFILLER_162_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6331_ _3069_ dmmu1.page_table\[3\]\[4\] _3077_ _3084_ vssd1 vssd1 vccd1 vccd1 _0500_
+ sky130_fd_sc_hd__a31o_1
XFILLER_162_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3543_ _0879_ _1122_ _1126_ _1127_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__a22o_1
XFILLER_127_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3815__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6262_ _2793_ _3040_ vssd1 vssd1 vccd1 vccd1 _3044_ sky130_fd_sc_hd__and2_1
XFILLER_282_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3474_ dmmu1.page_table\[12\]\[6\] dmmu1.page_table\[13\]\[6\] dmmu1.page_table\[14\]\[6\]
+ dmmu1.page_table\[15\]\[6\] _0858_ _0861_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__mux4_1
XANTENNA__7226__CLK clknet_leaf_22_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5213_ _2416_ dmmu0.page_table\[8\]\[9\] _2411_ vssd1 vssd1 vccd1 vccd1 _2422_ sky130_fd_sc_hd__and3_1
XFILLER_170_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6193_ _2879_ _3002_ vssd1 vssd1 vccd1 vccd1 _3003_ sky130_fd_sc_hd__and2_1
XFILLER_130_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5144_ _2371_ dmmu0.page_table\[10\]\[7\] _2373_ vssd1 vssd1 vccd1 vccd1 _2381_ sky130_fd_sc_hd__and3_1
XFILLER_130_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5075_ _2332_ immu_0.page_table\[12\]\[1\] _2336_ _2339_ vssd1 vssd1 vccd1 vccd1
+ _0798_ sky130_fd_sc_hd__a31o_1
XFILLER_151_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3619__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4026_ _1535_ _1536_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__and2_1
XFILLER_244_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6033__A1 _2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_18_core_clock_A clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5977_ _2867_ dmmu1.page_table\[13\]\[7\] _2859_ _2870_ vssd1 vssd1 vccd1 vccd1 _0360_
+ sky130_fd_sc_hd__a31o_1
XFILLER_197_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3398__A2 _0929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4928_ net94 vssd1 vssd1 vccd1 vccd1 _2251_ sky130_fd_sc_hd__buf_4
XANTENNA__4812__C _2174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4859_ _2182_ immu_1.page_table\[3\]\[3\] _2197_ vssd1 vssd1 vccd1 vccd1 _2201_ sky130_fd_sc_hd__and3_1
XFILLER_20_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6529_ clknet_leaf_41_core_clock _0599_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_118_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4320__S _1493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3858__A0 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4556__A _1981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6474__C _3159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input221_A dcache_mem_o_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input319_A ic0_wb_adr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6024__A1 _2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5387__A _1933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4291__A _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6893__CLK clknet_leaf_76_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4889__A2 _2219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6011__A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_20_core_clock_A clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_98_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output440_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output538_A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4510__A1 _1976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3190_ _0812_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__inv_6
XFILLER_182_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6263__A1 _3042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4813__A2 _2172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5900_ _1948_ _2812_ _2825_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__a21o_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6880_ clknet_leaf_70_core_clock _0141_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[5\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_201_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_9_core_clock_A clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5831_ _1950_ _2766_ _2781_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__a21o_1
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5369__A3 _2510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5762_ _2242_ _2730_ _2741_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__a21o_1
XANTENNA__4121__S0 _1493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7501_ net403 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_1
X_4713_ _2106_ immu_1.page_table\[9\]\[9\] _2103_ vssd1 vssd1 vccd1 vccd1 _2115_ sky130_fd_sc_hd__and3_1
XFILLER_187_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5693_ _2701_ vssd1 vssd1 vccd1 vccd1 _2702_ sky130_fd_sc_hd__buf_2
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4644_ _2010_ _2066_ _2073_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__a21o_1
X_7432_ net393 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_1
XFILLER_190_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5744__B _2572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4575_ _2029_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__clkbuf_4
X_7363_ net286 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_2
XFILLER_128_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6616__CLK clknet_leaf_54_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6314_ _3069_ dmmu1.page_table\[4\]\[11\] _3057_ _3073_ vssd1 vssd1 vccd1 vccd1 _0494_
+ sky130_fd_sc_hd__a31o_1
X_3526_ _1103_ _1104_ _1111_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__and3_1
X_7294_ clknet_leaf_43_core_clock _0555_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5829__A1 _1948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6245_ _3026_ dmmu1.page_table\[6\]\[9\] _3019_ _3032_ vssd1 vssd1 vccd1 vccd1 _0466_
+ sky130_fd_sc_hd__a31o_1
XFILLER_89_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3457_ dmmu0.page_table\[10\]\[5\] dmmu0.page_table\[11\]\[5\] _0910_ vssd1 vssd1
+ vccd1 vccd1 _1045_ sky130_fd_sc_hd__mux2_1
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6176_ _2977_ dmmu1.page_table\[8\]\[7\] _2981_ _2991_ vssd1 vssd1 vccd1 vccd1 _0438_
+ sky130_fd_sc_hd__a31o_1
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3388_ dmmu1.page_table\[12\]\[3\] dmmu1.page_table\[13\]\[3\] dmmu1.page_table\[14\]\[3\]
+ dmmu1.page_table\[15\]\[3\] _0892_ _0864_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__mux4_1
XFILLER_57_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5127_ _2370_ vssd1 vssd1 vccd1 vccd1 _2371_ sky130_fd_sc_hd__buf_2
XFILLER_257_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5058_ _2316_ immu_0.page_table\[14\]\[6\] _2320_ _2328_ vssd1 vssd1 vccd1 vccd1
+ _0792_ sky130_fd_sc_hd__a31o_1
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4009_ _1518_ _1519_ _1520_ _1447_ _1457_ vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__a221o_2
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6006__A1 _2884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4568__A1 _2023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4315__S _1493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4542__C _2004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5935__A _2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3455__A _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4050__S _1448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input171_A c1_o_req_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3543__A2 _1122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input269_A dcache_wb_o_dat[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6493__A1 _1979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput310 ic0_wb_adr[10] vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_1
XFILLER_283_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput321 ic0_wb_adr[6] vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input32_A c0_o_mem_data[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput332 ic1_mem_data[10] vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_86_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput343 ic1_mem_data[20] vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__buf_2
XFILLER_282_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput354 ic1_mem_data[30] vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_2
Xinput365 ic1_wb_adr[11] vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_2
XANTENNA__3190__A _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6245__A1 _3026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput376 ic1_wb_adr[7] vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput387 inner_wb_ack vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_8
XFILLER_208_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput398 inner_wb_i_dat[3] vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_8
XFILLER_275_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4559__A1 _2016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7071__CLK clknet_leaf_79_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5845__A _2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6639__CLK clknet_leaf_56_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5523__A3 _2607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4360_ _1857_ _1859_ _1861_ _1863_ _1457_ vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__a221o_2
XANTENNA__4192__C1 _1451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5283__C _2464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4731__A1 _2010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3311_ dmmu0.page_table\[4\]\[0\] dmmu0.page_table\[5\]\[0\] dmmu0.page_table\[6\]\[0\]
+ dmmu0.page_table\[7\]\[0\] _0900_ _0902_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__mux4_1
XFILLER_259_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4291_ _1430_ _1795_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__or2_1
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6030_ _2879_ _2904_ vssd1 vssd1 vccd1 vccd1 _2905_ sky130_fd_sc_hd__and2_1
X_3242_ net126 net21 _0840_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__mux2_1
XFILLER_86_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6395__B _3118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4798__A1 _2021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6932_ clknet_leaf_57_core_clock _0193_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_242_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6863_ clknet_leaf_71_core_clock _0124_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3470__A1 _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4135__S _1601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5814_ _2226_ _2767_ _2772_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__a21o_1
XFILLER_179_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6794_ clknet_leaf_10_core_clock _0055_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5745_ _2731_ vssd1 vssd1 vccd1 vccd1 _2732_ sky130_fd_sc_hd__buf_2
XANTENNA__5755__A _2736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4970__A1 _1972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4970__B2 immu_1.page_table\[0\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5676_ _1928_ immu_0.high_addr_off\[1\] _2690_ vssd1 vssd1 vccd1 vccd1 _2692_ sky130_fd_sc_hd__mux2_1
XFILLER_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5474__B _2577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7415_ net330 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__clkbuf_2
X_4627_ _2054_ immu_1.page_table\[12\]\[10\] _2048_ vssd1 vssd1 vccd1 vccd1 _2061_
+ sky130_fd_sc_hd__and3_1
XFILLER_190_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3275__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4558_ _2017_ immu_1.page_table\[14\]\[6\] _2004_ vssd1 vssd1 vccd1 vccd1 _2018_
+ sky130_fd_sc_hd__and3_1
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7346_ net288 vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_2
XFILLER_116_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3509_ _1093_ _1094_ _1034_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__o21ai_2
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4489_ net201 vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__buf_6
X_7277_ clknet_leaf_18_core_clock _0538_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5490__A _1929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6475__A1 _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5278__A2 _2462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6228_ _3010_ dmmu1.page_table\[6\]\[1\] _3019_ _3023_ vssd1 vssd1 vccd1 vccd1 _0458_
+ sky130_fd_sc_hd__a31o_1
XFILLER_89_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6159_ _1968_ _2978_ vssd1 vssd1 vccd1 vccd1 _2982_ sky130_fd_sc_hd__nor2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4789__A1 _2012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4834__A _1896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7094__CLK clknet_leaf_11_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3884__S _1390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4961__A1 _1989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input386_A inner_ext_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5384__B _2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput140 c1_o_mem_data[15] vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_2
XFILLER_236_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput151 c1_o_mem_high_addr[1] vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_209_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput162 c1_o_mem_we vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__buf_2
Xinput173 c1_o_req_addr[3] vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_1
Xinput184 c1_sr_bus_addr[12] vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_1
Xinput195 c1_sr_bus_addr[8] vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4744__A _2105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5559__B _2212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3452__A1 dmmu0.page_table\[1\]\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3860_ _1384_ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_1
XFILLER_189_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3791_ _1346_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4401__A0 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5575__A _2217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5530_ net100 _2609_ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__and2_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3807__B _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5461_ net83 net76 _2439_ vssd1 vssd1 vccd1 vccd1 _2572_ sky130_fd_sc_hd__or3_4
X_7200_ clknet_leaf_22_core_clock _0461_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4412_ net213 _0835_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__and2_1
XANTENNA__4704__A1 _2012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput603 net603 vssd1 vssd1 vccd1 vccd1 ic0_mem_ppl_submit sky130_fd_sc_hd__buf_2
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5392_ _1937_ _2527_ vssd1 vssd1 vccd1 vccd1 _2532_ sky130_fd_sc_hd__and2_1
Xoutput614 net614 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[15] sky130_fd_sc_hd__buf_2
XFILLER_132_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput625 net625 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[0] sky130_fd_sc_hd__buf_2
Xoutput636 net636 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[5] sky130_fd_sc_hd__buf_2
XFILLER_99_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput647 net647 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[0] sky130_fd_sc_hd__buf_2
XFILLER_259_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7131_ clknet_leaf_14_core_clock _0392_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4343_ immu_0.page_table\[4\]\[10\] immu_0.page_table\[5\]\[10\] _1472_ vssd1 vssd1
+ vccd1 vccd1 _1847_ sky130_fd_sc_hd__mux2_1
XFILLER_160_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput658 net658 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[5] sky130_fd_sc_hd__buf_2
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput669 net669 vssd1 vssd1 vccd1 vccd1 inner_wb_adr[13] sky130_fd_sc_hd__buf_2
XANTENNA__4919__A _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7062_ clknet_leaf_10_core_clock _0323_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4274_ _1462_ _1770_ _1779_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__or3b_1
XFILLER_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_274_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6013_ _2884_ dmmu1.page_table\[12\]\[8\] _2878_ _2892_ vssd1 vssd1 vccd1 vccd1 _0374_
+ sky130_fd_sc_hd__a31o_1
XFILLER_100_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3225_ _0833_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_1
XFILLER_140_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6209__A1 _3010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6915_ clknet_leaf_76_core_clock _0176_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3443__A1 _0869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6846_ clknet_leaf_69_core_clock _0107_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[8\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3994__A2 _1505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6954__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6777_ clknet_leaf_81_core_clock _0038_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3989_ immu_0.page_table\[2\]\[2\] immu_0.page_table\[3\]\[2\] _1472_ vssd1 vssd1
+ vccd1 vccd1 _1501_ sky130_fd_sc_hd__mux2_1
XANTENNA__5916__C _2832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5728_ immu_1.high_addr_off\[1\] _1967_ _2720_ vssd1 vssd1 vccd1 vccd1 _2722_ sky130_fd_sc_hd__mux2_1
XFILLER_210_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4820__C _2174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5659_ _2245_ _2669_ _2680_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__a21o_1
XFILLER_136_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4829__A _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5120__A1 _2363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3357__S1 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input134_A c1_o_mem_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3879__S _1386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4564__A _2017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input301_A ic0_mem_data[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__A2 _1477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3908__A _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4730__C _2123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3293__S0 _0865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6003__B _2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_core_clock clknet_3_4_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5842__B _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5111__A1 _2347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6827__CLK clknet_leaf_68_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6977__CLK clknet_leaf_11_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4961_ _1989_ _2256_ _2271_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__a21o_1
XANTENNA__3425__A1 _0918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6700_ clknet_leaf_42_core_clock _0770_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_189_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3912_ immu_0.page_table\[12\]\[0\] immu_0.page_table\[13\]\[0\] _1425_ vssd1 vssd1
+ vccd1 vccd1 _1426_ sky130_fd_sc_hd__mux2_1
X_4892_ _2204_ dmmu0.page_table\[0\]\[1\] _2221_ vssd1 vssd1 vccd1 vccd1 _2225_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_54_core_clock clknet_3_6_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5178__A1 _2243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6631_ clknet_leaf_55_core_clock _0701_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3843_ _1373_ net257 vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__and2_4
XFILLER_165_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6562_ clknet_leaf_49_core_clock _0632_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3774_ net161 net56 _0839_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__mux2_1
XANTENNA__4640__C _2068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6390__A3 _3116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5513_ _2561_ vssd1 vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__clkbuf_4
XFILLER_218_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6493_ dmmu1.long_off_reg\[5\] _1979_ _3172_ vssd1 vssd1 vccd1 vccd1 _3178_ sky130_fd_sc_hd__mux2_1
XFILLER_157_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5444_ _2562_ immu_0.page_table\[5\]\[2\] _2557_ _2563_ vssd1 vssd1 vccd1 vccd1 _0134_
+ sky130_fd_sc_hd__a31o_1
XFILLER_218_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput411 net411 vssd1 vssd1 vccd1 vccd1 c0_i_mem_ack sky130_fd_sc_hd__buf_2
XFILLER_145_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput422 net422 vssd1 vssd1 vccd1 vccd1 c0_i_mem_data[4] sky130_fd_sc_hd__buf_2
Xoutput433 net433 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[13] sky130_fd_sc_hd__buf_2
XFILLER_218_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput444 net444 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[23] sky130_fd_sc_hd__buf_2
XANTENNA__4649__A _2072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5375_ _2517_ immu_0.page_table\[8\]\[8\] _2510_ _2521_ vssd1 vssd1 vccd1 vccd1 _0107_
+ sky130_fd_sc_hd__a31o_1
Xoutput455 net455 vssd1 vssd1 vccd1 vccd1 c0_i_req_data[4] sky130_fd_sc_hd__buf_2
Xoutput466 net466 vssd1 vssd1 vccd1 vccd1 c1_i_core_int_sreg[1] sky130_fd_sc_hd__buf_2
X_7114_ clknet_leaf_31_core_clock _0375_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[12\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput477 net477 vssd1 vssd1 vccd1 vccd1 c1_i_mem_data[2] sky130_fd_sc_hd__buf_2
Xoutput488 net488 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[11] sky130_fd_sc_hd__buf_2
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4326_ _1569_ net244 _1805_ _1830_ vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__a22o_4
Xoutput499 net499 vssd1 vssd1 vccd1 vccd1 c1_i_req_data[21] sky130_fd_sc_hd__buf_2
XFILLER_86_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4257_ _1581_ _1762_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__nor2_1
X_7045_ clknet_leaf_36_core_clock _0306_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5653__A2 _2669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3208_ net224 _0824_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__and2_1
XFILLER_170_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4188_ _1581_ _1692_ _1694_ _1456_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__o211a_1
XFILLER_262_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3664__A1 _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_93_core_clock clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3416__A1 _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3511__S1 _0902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5169__A1 _2230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6829_ clknet_leaf_69_core_clock _0090_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4831__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7132__CLK clknet_leaf_34_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5646__C _2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3463__A _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3352__A0 _0864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_core_clock_A clknet_3_5_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_input251_A dcache_wb_adr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5892__A2 _2812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input349_A ic1_mem_data[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4447__A3 _1924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3655__A1 _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A2 _1468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5837__B _2278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4368__C1 _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6014__A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6372__A3 _3096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5580__A1 _2211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5853__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3490_ net46 dmmu0.long_off_reg\[1\] vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__xor2_1
XFILLER_185_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5160_ _2216_ _2388_ vssd1 vssd1 vccd1 vccd1 _2391_ sky130_fd_sc_hd__or2_1
XANTENNA__5883__A2 _2812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4111_ _1619_ vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__inv_2
XFILLER_284_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5091_ _2312_ _2338_ vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__and2_1
XFILLER_110_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4042_ net369 vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__buf_4
XANTENNA__4438__A3 _1924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7005__CLK clknet_leaf_36_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4843__B1 _2192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5399__A1 _2531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5993_ _2880_ vssd1 vssd1 vccd1 vccd1 _2881_ sky130_fd_sc_hd__buf_2
XFILLER_224_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7155__CLK clknet_leaf_30_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3949__A2 _1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4932__A _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4944_ _2262_ immu_1.page_table\[7\]\[2\] _2259_ vssd1 vssd1 vccd1 vccd1 _2263_ sky130_fd_sc_hd__and3_1
XFILLER_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4875_ _1989_ _2194_ _2209_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__a21o_1
XFILLER_32_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6614_ clknet_leaf_54_core_clock _0684_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[5\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3826_ _1363_ net264 vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__and2_1
XFILLER_165_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6545_ clknet_leaf_50_core_clock _0615_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5571__A1 _2242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3757_ _1328_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5763__A _2736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6476_ _2190_ immu_1.page_table\[8\]\[9\] _3159_ vssd1 vssd1 vccd1 vccd1 _3169_ sky130_fd_sc_hd__and3_1
X_3688_ _0859_ _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__or2_1
XFILLER_106_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5482__B _2577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4379__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5427_ _2310_ _2543_ vssd1 vssd1 vccd1 vccd1 _2552_ sky130_fd_sc_hd__and2_1
XANTENNA__5323__A1 _2489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4126__A2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3283__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5358_ _1930_ _2407_ vssd1 vssd1 vccd1 vccd1 _2512_ sky130_fd_sc_hd__nor2_4
XFILLER_87_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3885__A1 _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4309_ _1496_ _1811_ _1813_ _1516_ vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__o211a_1
XFILLER_275_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5289_ _2458_ dmmu0.page_table\[14\]\[7\] _2464_ vssd1 vssd1 vccd1 vccd1 _2472_ sky130_fd_sc_hd__and3_1
XANTENNA__5626__A2 _2650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7028_ clknet_leaf_82_core_clock _0289_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[13\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_261_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4318__S _1493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5003__A _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4545__C _2004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6522__CLK clknet_leaf_43_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input299_A ic0_mem_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6672__CLK clknet_leaf_58_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3573__B1 _0872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6106__A3 _2942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5392__B _2527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input62_A c0_o_req_addr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5314__A1 _2363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3193__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7028__CLK clknet_leaf_82_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3876__A1 _1395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3971__S1 _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7178__CLK clknet_leaf_33_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_253_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6009__A _2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5848__A _2793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4752__A _2134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3487__S0 _0900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4471__B _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_core_clock clknet_3_1_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4660_ _2000_ _2081_ vssd1 vssd1 vccd1 vccd1 _2082_ sky130_fd_sc_hd__nor2_1
XFILLER_187_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_93_core_clock_A clknet_3_0_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3611_ _0993_ _1168_ _1194_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__o21a_4
XANTENNA__5553__A1 _2235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4591_ _2038_ immu_1.page_table\[13\]\[6\] _2032_ vssd1 vssd1 vccd1 vccd1 _2040_
+ sky130_fd_sc_hd__and3_1
XANTENNA__5583__A _2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3564__B1 _0872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6330_ net204 _3079_ vssd1 vssd1 vccd1 vccd1 _3084_ sky130_fd_sc_hd__and2_1
X_3542_ _1123_ _1124_ _1125_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__a21o_1
XFILLER_127_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3815__B _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5305__A1 _2363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6261_ _3042_ dmmu1.page_table\[5\]\[1\] _3038_ _3043_ vssd1 vssd1 vccd1 vccd1 _0471_
+ sky130_fd_sc_hd__a31o_1
X_3473_ _1058_ _1059_ _0881_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__mux2_1
XFILLER_182_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5212_ _2245_ _2409_ _2421_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__a21o_1
XFILLER_142_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6192_ _3001_ vssd1 vssd1 vccd1 vccd1 _3002_ sky130_fd_sc_hd__clkbuf_4
XFILLER_269_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5143_ _2240_ _2369_ _2380_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__a21o_1
XFILLER_111_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5074_ _1928_ _2338_ vssd1 vssd1 vccd1 vccd1 _2339_ sky130_fd_sc_hd__and2_1
XFILLER_84_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3619__A1 _0868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4025_ immu_0.page_table\[8\]\[3\] immu_0.page_table\[9\]\[3\] immu_0.page_table\[10\]\[3\]
+ immu_0.page_table\[11\]\[3\] _1472_ _1419_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__mux4_1
XFILLER_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6545__CLK clknet_leaf_50_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3977__S _1443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4662__A _1998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5976_ _2803_ _2861_ vssd1 vssd1 vccd1 vccd1 _2870_ sky130_fd_sc_hd__and2_1
XFILLER_40_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4927_ _2249_ _2218_ _2250_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__a21o_1
XFILLER_200_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3278__A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6695__CLK clknet_leaf_42_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5196__C _2411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4858_ _1972_ _2195_ _2200_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__a21o_1
XANTENNA__6336__A3 _3077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3809_ net218 _1348_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__and2_1
X_4789_ _2012_ _2155_ _2162_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__a21o_1
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6528_ clknet_leaf_41_core_clock _0598_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5924__C _2832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6459_ _1995_ _3157_ _3160_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__a21o_1
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5075__A3 _2336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input214_A dcache_mem_o_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3887__S _1390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5668__A _2682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4572__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4035__A1 _1419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5387__B _2527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5783__A1 _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3188__A _0811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6327__A3 _3077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5535__A1 _2603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6499__A _1914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3916__A _1419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output433_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6568__CLK clknet_leaf_49_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5830_ _2777_ dmmu0.page_table\[3\]\[10\] _2768_ vssd1 vssd1 vccd1 vccd1 _2781_ sky130_fd_sc_hd__and3_1
XFILLER_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4913__C _2221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5761_ _2736_ dmmu0.page_table\[4\]\[7\] _2732_ vssd1 vssd1 vccd1 vccd1 _2741_ sky130_fd_sc_hd__and3_1
XANTENNA__4121__S1 _1442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7500_ net402 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_1
X_4712_ _2021_ _2101_ _2114_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__a21o_1
XFILLER_277_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5692_ _2443_ _2605_ vssd1 vssd1 vccd1 vccd1 _2701_ sky130_fd_sc_hd__or2_1
XFILLER_202_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7431_ net392 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_1
X_4643_ _2072_ immu_1.page_table\[11\]\[3\] _2068_ vssd1 vssd1 vccd1 vccd1 _2073_
+ sky130_fd_sc_hd__and3_1
XANTENNA__3826__A _1363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7362_ net285 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_2
X_4574_ _2000_ _2028_ vssd1 vssd1 vccd1 vccd1 _2029_ sky130_fd_sc_hd__nor2_1
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6313_ net199 _3059_ vssd1 vssd1 vccd1 vccd1 _3073_ sky130_fd_sc_hd__and2_1
XFILLER_190_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3525_ _1109_ _1110_ _0957_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__o21ai_1
X_7293_ clknet_leaf_43_core_clock _0554_ vssd1 vssd1 vccd1 vccd1 immu_1.page_table\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6244_ _2893_ _3021_ vssd1 vssd1 vccd1 vccd1 _3032_ sky130_fd_sc_hd__and2_1
XFILLER_143_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3456_ _0918_ _1041_ _1043_ _0899_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__a31o_1
XFILLER_170_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4657__A _2072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6175_ _2803_ _2983_ vssd1 vssd1 vccd1 vccd1 _2991_ sky130_fd_sc_hd__and2_1
X_3387_ dmmu1.page_table\[8\]\[3\] dmmu1.page_table\[9\]\[3\] dmmu1.page_table\[10\]\[3\]
+ dmmu1.page_table\[11\]\[3\] _0892_ _0864_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__mux4_1
XANTENNA__3561__A _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5126_ _1896_ vssd1 vssd1 vccd1 vccd1 _2370_ sky130_fd_sc_hd__buf_2
XFILLER_84_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5057_ _1942_ _2322_ vssd1 vssd1 vccd1 vccd1 _2328_ sky130_fd_sc_hd__and2_1
XFILLER_284_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4008_ immu_1.page_table\[8\]\[2\] immu_1.page_table\[9\]\[2\] _1443_ vssd1 vssd1
+ vccd1 vccd1 _1520_ sky130_fd_sc_hd__mux2_1
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5488__A _2561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4823__C _2174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4568__A2 _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5959_ _1968_ _2028_ vssd1 vssd1 vccd1 vccd1 _2860_ sky130_fd_sc_hd__nor2_1
XFILLER_80_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5654__C _2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input164_A c1_o_req_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6710__CLK clknet_leaf_63_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4567__A _2017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput300 ic0_mem_data[30] vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_1
XFILLER_248_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput311 ic0_wb_adr[11] vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_1
XFILLER_96_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput322 ic0_wb_adr[7] vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_2
Xinput333 ic1_mem_data[11] vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_2
XFILLER_29_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input331_A ic1_mem_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput344 ic1_mem_data[21] vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_2
XFILLER_48_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput355 ic1_mem_data[31] vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_2
XFILLER_236_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput366 ic1_wb_adr[12] vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__buf_2
Xinput377 ic1_wb_adr[8] vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_2
XANTENNA__5048__A3 _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input25_A c0_o_mem_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput388 inner_wb_err vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_8
Xinput399 inner_wb_i_dat[4] vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_8
XANTENNA__6860__CLK clknet_leaf_71_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3464__C1 _0906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5398__A _1944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7216__CLK clknet_leaf_22_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4559__A2 _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5756__A1 _2232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5845__B _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5508__A1 _2588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6022__A _2561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4731__A2 _2120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3310_ dmmu0.page_table\[0\]\[0\] dmmu0.page_table\[1\]\[0\] dmmu0.page_table\[2\]\[0\]
+ dmmu0.page_table\[3\]\[0\] _0900_ _0902_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__mux4_1
XFILLER_125_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4290_ immu_0.page_table\[8\]\[9\] immu_0.page_table\[9\]\[9\] _1425_ vssd1 vssd1
+ vccd1 vccd1 _1795_ sky130_fd_sc_hd__mux2_1
XFILLER_152_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3241_ _0843_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_258_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4247__A1 _1479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6931_ clknet_leaf_77_core_clock _0192_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_214_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5995__A1 _2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4798__A2 _2155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_2_1_core_clock clknet_opt_2_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_opt_2_1_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6862_ clknet_leaf_70_core_clock _0123_ vssd1 vssd1 vccd1 vccd1 immu_0.page_table\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4643__C _2068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5101__A _1930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3470__A2 _1035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5813_ _2762_ dmmu0.page_table\[3\]\[2\] _2769_ vssd1 vssd1 vccd1 vccd1 _2772_ sky130_fd_sc_hd__and3_1
XFILLER_222_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5747__A1 _2210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6793_ clknet_leaf_80_core_clock _0054_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3758__A0 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5744_ _2443_ _2572_ vssd1 vssd1 vccd1 vccd1 _2731_ sky130_fd_sc_hd__or2_1
XFILLER_210_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5675_ _2691_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4970__A2 _2274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7414_ net355 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4151__S _1453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4626_ _2023_ _2047_ _2060_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__a21o_1
XFILLER_135_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6172__A1 _2977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6733__CLK clknet_leaf_63_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7345_ net277 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_2
X_4557_ _1897_ vssd1 vssd1 vccd1 vccd1 _2017_ sky130_fd_sc_hd__clkbuf_4
XFILLER_150_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5771__A _2736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3508_ _1089_ _1090_ _1092_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__and3_1
X_7276_ clknet_leaf_22_core_clock _0537_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4488_ _1939_ dmmu1.page_table\[14\]\[0\] _1964_ _1966_ vssd1 vssd1 vccd1 vccd1 _0584_
+ sky130_fd_sc_hd__a31o_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5490__B _2589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6475__A2 _3157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6227_ _2791_ _3021_ vssd1 vssd1 vccd1 vccd1 _3023_ sky130_fd_sc_hd__and2_1
XFILLER_77_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3439_ dmmu1.page_table\[8\]\[5\] dmmu1.page_table\[9\]\[5\] dmmu1.page_table\[10\]\[5\]
+ dmmu1.page_table\[11\]\[5\] _0892_ _0864_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__mux4_1
XFILLER_277_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4818__C _2174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6158_ _2980_ vssd1 vssd1 vccd1 vccd1 _2981_ sky130_fd_sc_hd__clkbuf_4
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3694__C1 _0854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5109_ _2347_ immu_0.page_table\[13\]\[4\] _2353_ _2359_ vssd1 vssd1 vccd1 vccd1
+ _0003_ sky130_fd_sc_hd__a31o_1
XFILLER_57_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6089_ _1993_ _2923_ vssd1 vssd1 vccd1 vccd1 _2939_ sky130_fd_sc_hd__and2_1
XFILLER_272_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4238__A1 _1570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4789__A2 _2155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5450__A3 _2557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6107__A _2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5011__A _1926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5738__A1 _1981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4097__S0 _1601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input281_A ic0_mem_data[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input379_A ic1_wb_cyc vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4174__B1 _1654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1_0_core_clock clknet_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_1_1_0_core_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_107_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5674__A0 _2210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4728__C _2123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput130 c1_o_mem_addr[6] vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
XFILLER_76_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput141 c1_o_mem_data[1] vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_2
XFILLER_248_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput152 c1_o_mem_high_addr[2] vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput163 c1_o_req_active vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
XFILLER_248_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput174 c1_o_req_addr[4] vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_1
Xinput185 c1_sr_bus_addr[13] vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_1
XANTENNA__7401__A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput196 c1_sr_bus_addr[9] vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5977__A1 _2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3437__C1 _0855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4236__S _1408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6606__CLK clknet_leaf_62_core_clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6017__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_core_clock clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_core_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_32_core_clock_A clknet_3_7_0_core_clock vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4760__A _2134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3790_ net224 _0993_ vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__and2_1
XANTENNA__4401__A1 _1899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5575__B _2334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5294__C _2464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5460_ _2562_ immu_0.page_table\[5\]\[10\] _2556_ _2571_ vssd1 vssd1 vccd1 vccd1
+ _0142_ sky130_fd_sc_hd__a31o_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4411_ _1905_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_2
XANTENNA__4704__A2 _2101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput604 net604 vssd1 vssd1 vccd1 vccd1 ic0_mem_req sky130_fd_sc_hd__buf_2
XFILLER_172_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput615 net615 vssd1 vssd1 vccd1 vccd1 ic0_wb_i_dat[1] sky130_fd_sc_hd__buf_2
X_5391_ _2300_ vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__clkbuf_4
Xoutput626 net626 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[10] sky130_fd_sc_hd__buf_2
XFILLER_160_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7130_ clknet_leaf_29_core_clock _0391_ vssd1 vssd1 vccd1 vccd1 dmmu1.page_table\[11\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput637 net637 vssd1 vssd1 vccd1 vccd1 ic1_mem_addr[6] sky130_fd_sc_hd__buf_2
Xoutput648 net648 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[10] sky130_fd_sc_hd__buf_2
X_4342_ _1424_ _1845_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__or2_1
XFILLER_113_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput659 net659 vssd1 vssd1 vccd1 vccd1 ic1_wb_i_dat[6] sky130_fd_sc_hd__buf_2
XFILLER_125_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7061_ clknet_leaf_80_core_clock _0322_ vssd1 vssd1 vccd1 vccd1 dmmu0.page_table\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4273_ _1516_ _1772_ _1774_ _1778_ _1553_ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__a311o_1
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4638__C _2068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6012_ _2891_ _2881_ vssd1 vssd1 vccd1 vccd1 _2892_ sky130_fd_sc_hd__and2_1
XFILLER_39_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4000__A _1419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3224_ net217 _0824_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__and2_1
.ends

