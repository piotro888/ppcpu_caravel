module interconnect_outer (c0_clk,
    c1_clk,
    dcache_clk,
    ic0_clk,
    ic1_clk,
    inner_clock,
    inner_disable,
    inner_embed_mode,
    inner_ext_irq,
    inner_reset,
    inner_wb_4_burst,
    inner_wb_8_burst,
    inner_wb_ack,
    inner_wb_cyc,
    inner_wb_err,
    inner_wb_stb,
    inner_wb_we,
    iram_clk,
    iram_we,
    mgt_wb_ack_o,
    mgt_wb_clk_i,
    mgt_wb_cyc_i,
    mgt_wb_rst_i,
    mgt_wb_stb_i,
    mgt_wb_we_i,
    user_clock2,
    vccd1,
    vssd1,
    inner_wb_adr,
    inner_wb_i_dat,
    inner_wb_o_dat,
    inner_wb_sel,
    iram_addr,
    iram_i_data,
    iram_o_data,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    m_io_in,
    m_io_oeb,
    m_io_out,
    mgt_wb_adr_i,
    mgt_wb_dat_i,
    mgt_wb_dat_o,
    mgt_wb_sel_i);
 output c0_clk;
 output c1_clk;
 output dcache_clk;
 output ic0_clk;
 output ic1_clk;
 output inner_clock;
 output inner_disable;
 output inner_embed_mode;
 output inner_ext_irq;
 output inner_reset;
 input inner_wb_4_burst;
 input inner_wb_8_burst;
 output inner_wb_ack;
 input inner_wb_cyc;
 output inner_wb_err;
 input inner_wb_stb;
 input inner_wb_we;
 output iram_clk;
 output iram_we;
 output mgt_wb_ack_o;
 input mgt_wb_clk_i;
 input mgt_wb_cyc_i;
 input mgt_wb_rst_i;
 input mgt_wb_stb_i;
 input mgt_wb_we_i;
 input user_clock2;
 input vccd1;
 input vssd1;
 input [23:0] inner_wb_adr;
 output [15:0] inner_wb_i_dat;
 input [15:0] inner_wb_o_dat;
 input [1:0] inner_wb_sel;
 output [5:0] iram_addr;
 output [15:0] iram_i_data;
 input [15:0] iram_o_data;
 output [2:0] irq;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 input [37:0] m_io_in;
 output [37:0] m_io_oeb;
 output [37:0] m_io_out;
 input [31:0] mgt_wb_adr_i;
 input [31:0] mgt_wb_dat_i;
 output [31:0] mgt_wb_dat_o;
 input [3:0] mgt_wb_sel_i;

 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net269;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net270;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net271;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net272;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net273;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net379;
 wire net380;
 wire net334;
 wire net335;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net336;
 wire net337;
 wire net332;
 wire net333;
 wire net338;
 wire net339;
 wire net387;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net348;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net349;
 wire net377;
 wire net378;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire \clk_div.clock_sel ;
 wire \clk_div.clock_sel_r ;
 wire \clk_div.cnt[0] ;
 wire \clk_div.cnt[10] ;
 wire \clk_div.cnt[11] ;
 wire \clk_div.cnt[12] ;
 wire \clk_div.cnt[13] ;
 wire \clk_div.cnt[14] ;
 wire \clk_div.cnt[15] ;
 wire \clk_div.cnt[1] ;
 wire \clk_div.cnt[2] ;
 wire \clk_div.cnt[3] ;
 wire \clk_div.cnt[4] ;
 wire \clk_div.cnt[5] ;
 wire \clk_div.cnt[6] ;
 wire \clk_div.cnt[7] ;
 wire \clk_div.cnt[8] ;
 wire \clk_div.cnt[9] ;
 wire \clk_div.curr_div[0] ;
 wire \clk_div.curr_div[1] ;
 wire \clk_div.curr_div[2] ;
 wire \clk_div.curr_div[3] ;
 wire \clk_div.next_div_buff[0] ;
 wire \clk_div.next_div_buff[1] ;
 wire \clk_div.next_div_buff[2] ;
 wire \clk_div.next_div_buff[3] ;
 wire \clk_div.next_div_val ;
 wire \clk_div.res_clk ;
 wire clknet_0_net196;
 wire clknet_0_user_clock2;
 wire clknet_2_0__leaf_user_clock2;
 wire clknet_2_1__leaf_user_clock2;
 wire clknet_2_2__leaf_user_clock2;
 wire clknet_2_3__leaf_user_clock2;
 wire clknet_4_0_0_net196;
 wire clknet_4_10_0_net196;
 wire clknet_4_11_0_net196;
 wire clknet_4_12_0_net196;
 wire clknet_4_13_0_net196;
 wire clknet_4_14_0_net196;
 wire clknet_4_15_0_net196;
 wire clknet_4_1_0_net196;
 wire clknet_4_2_0_net196;
 wire clknet_4_3_0_net196;
 wire clknet_4_4_0_net196;
 wire clknet_4_5_0_net196;
 wire clknet_4_6_0_net196;
 wire clknet_4_7_0_net196;
 wire clknet_4_8_0_net196;
 wire clknet_4_9_0_net196;
 wire clknet_leaf_0_user_clock2;
 wire clknet_leaf_10_user_clock2;
 wire clknet_leaf_11_user_clock2;
 wire clknet_leaf_12_user_clock2;
 wire clknet_leaf_13_user_clock2;
 wire clknet_leaf_14_user_clock2;
 wire clknet_leaf_15_user_clock2;
 wire clknet_leaf_16_user_clock2;
 wire clknet_leaf_17_user_clock2;
 wire clknet_leaf_18_user_clock2;
 wire clknet_leaf_19_user_clock2;
 wire clknet_leaf_1_user_clock2;
 wire clknet_leaf_20_user_clock2;
 wire clknet_leaf_21_user_clock2;
 wire clknet_leaf_22_user_clock2;
 wire clknet_leaf_23_user_clock2;
 wire clknet_leaf_24_user_clock2;
 wire clknet_leaf_25_user_clock2;
 wire clknet_leaf_26_user_clock2;
 wire clknet_leaf_27_user_clock2;
 wire clknet_leaf_28_user_clock2;
 wire clknet_leaf_29_user_clock2;
 wire clknet_leaf_2_user_clock2;
 wire clknet_leaf_30_user_clock2;
 wire clknet_leaf_31_user_clock2;
 wire clknet_leaf_32_user_clock2;
 wire clknet_leaf_33_user_clock2;
 wire clknet_leaf_35_user_clock2;
 wire clknet_leaf_36_user_clock2;
 wire clknet_leaf_37_user_clock2;
 wire clknet_leaf_38_user_clock2;
 wire clknet_leaf_39_user_clock2;
 wire clknet_leaf_3_user_clock2;
 wire clknet_leaf_40_user_clock2;
 wire clknet_leaf_41_user_clock2;
 wire clknet_leaf_42_user_clock2;
 wire clknet_leaf_43_user_clock2;
 wire clknet_leaf_44_user_clock2;
 wire clknet_leaf_45_user_clock2;
 wire clknet_leaf_46_user_clock2;
 wire clknet_leaf_47_user_clock2;
 wire clknet_leaf_49_user_clock2;
 wire clknet_leaf_4_user_clock2;
 wire clknet_leaf_50_user_clock2;
 wire clknet_leaf_5_user_clock2;
 wire clknet_leaf_6_user_clock2;
 wire clknet_leaf_7_user_clock2;
 wire clknet_leaf_8_user_clock2;
 wire clknet_leaf_9_user_clock2;
 wire \disable_s_ff[0] ;
 wire \embed_s_ff[0] ;
 wire \iram_latched[0] ;
 wire \iram_latched[10] ;
 wire \iram_latched[11] ;
 wire \iram_latched[12] ;
 wire \iram_latched[13] ;
 wire \iram_latched[14] ;
 wire \iram_latched[15] ;
 wire \iram_latched[1] ;
 wire \iram_latched[2] ;
 wire \iram_latched[3] ;
 wire \iram_latched[4] ;
 wire \iram_latched[5] ;
 wire \iram_latched[6] ;
 wire \iram_latched[7] ;
 wire \iram_latched[8] ;
 wire \iram_latched[9] ;
 wire iram_wb_ack;
 wire iram_wb_ack_del;
 wire \irq_s_ff[0] ;
 wire \m_arbiter.i_wb0_cyc ;
 wire \m_arbiter.o_sel_sig ;
 wire \m_arbiter.wb0_adr[0] ;
 wire \m_arbiter.wb0_adr[10] ;
 wire \m_arbiter.wb0_adr[11] ;
 wire \m_arbiter.wb0_adr[12] ;
 wire \m_arbiter.wb0_adr[13] ;
 wire \m_arbiter.wb0_adr[14] ;
 wire \m_arbiter.wb0_adr[15] ;
 wire \m_arbiter.wb0_adr[16] ;
 wire \m_arbiter.wb0_adr[17] ;
 wire \m_arbiter.wb0_adr[18] ;
 wire \m_arbiter.wb0_adr[19] ;
 wire \m_arbiter.wb0_adr[1] ;
 wire \m_arbiter.wb0_adr[20] ;
 wire \m_arbiter.wb0_adr[21] ;
 wire \m_arbiter.wb0_adr[22] ;
 wire \m_arbiter.wb0_adr[23] ;
 wire \m_arbiter.wb0_adr[2] ;
 wire \m_arbiter.wb0_adr[3] ;
 wire \m_arbiter.wb0_adr[4] ;
 wire \m_arbiter.wb0_adr[5] ;
 wire \m_arbiter.wb0_adr[6] ;
 wire \m_arbiter.wb0_adr[7] ;
 wire \m_arbiter.wb0_adr[8] ;
 wire \m_arbiter.wb0_adr[9] ;
 wire \m_arbiter.wb0_o_dat[0] ;
 wire \m_arbiter.wb0_o_dat[10] ;
 wire \m_arbiter.wb0_o_dat[11] ;
 wire \m_arbiter.wb0_o_dat[12] ;
 wire \m_arbiter.wb0_o_dat[13] ;
 wire \m_arbiter.wb0_o_dat[14] ;
 wire \m_arbiter.wb0_o_dat[15] ;
 wire \m_arbiter.wb0_o_dat[1] ;
 wire \m_arbiter.wb0_o_dat[2] ;
 wire \m_arbiter.wb0_o_dat[3] ;
 wire \m_arbiter.wb0_o_dat[4] ;
 wire \m_arbiter.wb0_o_dat[5] ;
 wire \m_arbiter.wb0_o_dat[6] ;
 wire \m_arbiter.wb0_o_dat[7] ;
 wire \m_arbiter.wb0_o_dat[8] ;
 wire \m_arbiter.wb0_o_dat[9] ;
 wire \m_arbiter.wb0_we ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \rst_cw_sync.reset_sync_ff[0] ;
 wire \rst_cw_sync.reset_sync_ff[1] ;
 wire \rst_cw_sync.reset_sync_ff[2] ;
 wire \rst_soc_sync.reset_sync_ff[0] ;
 wire \rst_soc_sync.reset_sync_ff[1] ;
 wire \rst_soc_sync.reset_sync_ff[2] ;
 wire \split_s_ff[0] ;
 wire \sspi.bit_cnt[0] ;
 wire \sspi.bit_cnt[1] ;
 wire \sspi.bit_cnt[2] ;
 wire \sspi.bit_cnt[3] ;
 wire \sspi.bit_cnt[4] ;
 wire \sspi.req_addr[0] ;
 wire \sspi.req_addr[10] ;
 wire \sspi.req_addr[11] ;
 wire \sspi.req_addr[12] ;
 wire \sspi.req_addr[13] ;
 wire \sspi.req_addr[14] ;
 wire \sspi.req_addr[15] ;
 wire \sspi.req_addr[16] ;
 wire \sspi.req_addr[17] ;
 wire \sspi.req_addr[18] ;
 wire \sspi.req_addr[19] ;
 wire \sspi.req_addr[1] ;
 wire \sspi.req_addr[20] ;
 wire \sspi.req_addr[21] ;
 wire \sspi.req_addr[22] ;
 wire \sspi.req_addr[23] ;
 wire \sspi.req_addr[2] ;
 wire \sspi.req_addr[3] ;
 wire \sspi.req_addr[4] ;
 wire \sspi.req_addr[5] ;
 wire \sspi.req_addr[6] ;
 wire \sspi.req_addr[7] ;
 wire \sspi.req_addr[8] ;
 wire \sspi.req_addr[9] ;
 wire \sspi.req_data[0] ;
 wire \sspi.req_data[10] ;
 wire \sspi.req_data[11] ;
 wire \sspi.req_data[12] ;
 wire \sspi.req_data[13] ;
 wire \sspi.req_data[14] ;
 wire \sspi.req_data[15] ;
 wire \sspi.req_data[1] ;
 wire \sspi.req_data[2] ;
 wire \sspi.req_data[3] ;
 wire \sspi.req_data[4] ;
 wire \sspi.req_data[5] ;
 wire \sspi.req_data[6] ;
 wire \sspi.req_data[7] ;
 wire \sspi.req_data[8] ;
 wire \sspi.req_data[9] ;
 wire \sspi.res_data[0] ;
 wire \sspi.res_data[10] ;
 wire \sspi.res_data[11] ;
 wire \sspi.res_data[12] ;
 wire \sspi.res_data[13] ;
 wire \sspi.res_data[14] ;
 wire \sspi.res_data[15] ;
 wire \sspi.res_data[1] ;
 wire \sspi.res_data[2] ;
 wire \sspi.res_data[3] ;
 wire \sspi.res_data[4] ;
 wire \sspi.res_data[5] ;
 wire \sspi.res_data[6] ;
 wire \sspi.res_data[7] ;
 wire \sspi.res_data[8] ;
 wire \sspi.res_data[9] ;
 wire \sspi.resp_err ;
 wire \sspi.state[0] ;
 wire \sspi.state[1] ;
 wire \sspi.state[2] ;
 wire \sspi.state[3] ;
 wire \sspi.state[4] ;
 wire \sspi.state[5] ;
 wire \sspi.state[6] ;
 wire \sspi.state[7] ;
 wire \sspi.sy_clk[0] ;
 wire \sspi.sy_clk[1] ;
 wire \sspi.sy_clk[2] ;
 wire \sspi.sy_clk[3] ;
 wire \wb_compressor.burst_cnt[0] ;
 wire \wb_compressor.burst_cnt[1] ;
 wire \wb_compressor.burst_cnt[2] ;
 wire \wb_compressor.burst_end[0] ;
 wire \wb_compressor.burst_end[2] ;
 wire \wb_compressor.l_we ;
 wire \wb_compressor.state[0] ;
 wire \wb_compressor.state[1] ;
 wire \wb_compressor.state[2] ;
 wire \wb_compressor.state[3] ;
 wire \wb_compressor.state[4] ;
 wire \wb_compressor.state[5] ;
 wire \wb_compressor.state[6] ;
 wire \wb_compressor.wb_ack ;
 wire \wb_compressor.wb_err ;
 wire \wb_compressor.wb_i_dat[0] ;
 wire \wb_compressor.wb_i_dat[10] ;
 wire \wb_compressor.wb_i_dat[11] ;
 wire \wb_compressor.wb_i_dat[12] ;
 wire \wb_compressor.wb_i_dat[13] ;
 wire \wb_compressor.wb_i_dat[14] ;
 wire \wb_compressor.wb_i_dat[15] ;
 wire \wb_compressor.wb_i_dat[1] ;
 wire \wb_compressor.wb_i_dat[2] ;
 wire \wb_compressor.wb_i_dat[3] ;
 wire \wb_compressor.wb_i_dat[4] ;
 wire \wb_compressor.wb_i_dat[5] ;
 wire \wb_compressor.wb_i_dat[6] ;
 wire \wb_compressor.wb_i_dat[7] ;
 wire \wb_compressor.wb_i_dat[8] ;
 wire \wb_compressor.wb_i_dat[9] ;
 wire \wb_cross_clk.ack_next_hold ;
 wire \wb_cross_clk.ack_xor_flag ;
 wire \wb_cross_clk.err_xor_flag ;
 wire \wb_cross_clk.m_burst_cnt[0] ;
 wire \wb_cross_clk.m_burst_cnt[1] ;
 wire \wb_cross_clk.m_burst_cnt[2] ;
 wire \wb_cross_clk.m_burst_cnt[3] ;
 wire \wb_cross_clk.m_new_req_flag ;
 wire \wb_cross_clk.m_s_sync.d_data[0] ;
 wire \wb_cross_clk.m_s_sync.d_data[10] ;
 wire \wb_cross_clk.m_s_sync.d_data[11] ;
 wire \wb_cross_clk.m_s_sync.d_data[12] ;
 wire \wb_cross_clk.m_s_sync.d_data[13] ;
 wire \wb_cross_clk.m_s_sync.d_data[14] ;
 wire \wb_cross_clk.m_s_sync.d_data[15] ;
 wire \wb_cross_clk.m_s_sync.d_data[16] ;
 wire \wb_cross_clk.m_s_sync.d_data[17] ;
 wire \wb_cross_clk.m_s_sync.d_data[18] ;
 wire \wb_cross_clk.m_s_sync.d_data[19] ;
 wire \wb_cross_clk.m_s_sync.d_data[1] ;
 wire \wb_cross_clk.m_s_sync.d_data[20] ;
 wire \wb_cross_clk.m_s_sync.d_data[21] ;
 wire \wb_cross_clk.m_s_sync.d_data[22] ;
 wire \wb_cross_clk.m_s_sync.d_data[23] ;
 wire \wb_cross_clk.m_s_sync.d_data[24] ;
 wire \wb_cross_clk.m_s_sync.d_data[25] ;
 wire \wb_cross_clk.m_s_sync.d_data[26] ;
 wire \wb_cross_clk.m_s_sync.d_data[27] ;
 wire \wb_cross_clk.m_s_sync.d_data[28] ;
 wire \wb_cross_clk.m_s_sync.d_data[29] ;
 wire \wb_cross_clk.m_s_sync.d_data[2] ;
 wire \wb_cross_clk.m_s_sync.d_data[30] ;
 wire \wb_cross_clk.m_s_sync.d_data[31] ;
 wire \wb_cross_clk.m_s_sync.d_data[32] ;
 wire \wb_cross_clk.m_s_sync.d_data[33] ;
 wire \wb_cross_clk.m_s_sync.d_data[34] ;
 wire \wb_cross_clk.m_s_sync.d_data[35] ;
 wire \wb_cross_clk.m_s_sync.d_data[36] ;
 wire \wb_cross_clk.m_s_sync.d_data[37] ;
 wire \wb_cross_clk.m_s_sync.d_data[38] ;
 wire \wb_cross_clk.m_s_sync.d_data[39] ;
 wire \wb_cross_clk.m_s_sync.d_data[3] ;
 wire \wb_cross_clk.m_s_sync.d_data[40] ;
 wire \wb_cross_clk.m_s_sync.d_data[41] ;
 wire \wb_cross_clk.m_s_sync.d_data[42] ;
 wire \wb_cross_clk.m_s_sync.d_data[43] ;
 wire \wb_cross_clk.m_s_sync.d_data[44] ;
 wire \wb_cross_clk.m_s_sync.d_data[45] ;
 wire \wb_cross_clk.m_s_sync.d_data[46] ;
 wire \wb_cross_clk.m_s_sync.d_data[4] ;
 wire \wb_cross_clk.m_s_sync.d_data[5] ;
 wire \wb_cross_clk.m_s_sync.d_data[6] ;
 wire \wb_cross_clk.m_s_sync.d_data[7] ;
 wire \wb_cross_clk.m_s_sync.d_data[8] ;
 wire \wb_cross_clk.m_s_sync.d_data[9] ;
 wire \wb_cross_clk.m_s_sync.d_xfer_xor_sync[0] ;
 wire \wb_cross_clk.m_s_sync.d_xfer_xor_sync[1] ;
 wire \wb_cross_clk.m_s_sync.d_xfer_xor_sync[2] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[0] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[10] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[11] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[12] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[13] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[14] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[15] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[16] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[17] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[18] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[19] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[1] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[20] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[21] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[22] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[23] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[24] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[25] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[26] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[27] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[28] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[29] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[2] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[30] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[31] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[32] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[33] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[34] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[35] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[36] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[37] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[38] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[39] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[3] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[40] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[41] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[42] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[43] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[44] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[45] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[46] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[4] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[5] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[6] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[7] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[8] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[9] ;
 wire \wb_cross_clk.m_s_sync.s_xfer_xor_flag ;
 wire \wb_cross_clk.m_wb_i_dat[0] ;
 wire \wb_cross_clk.m_wb_i_dat[10] ;
 wire \wb_cross_clk.m_wb_i_dat[11] ;
 wire \wb_cross_clk.m_wb_i_dat[12] ;
 wire \wb_cross_clk.m_wb_i_dat[13] ;
 wire \wb_cross_clk.m_wb_i_dat[14] ;
 wire \wb_cross_clk.m_wb_i_dat[15] ;
 wire \wb_cross_clk.m_wb_i_dat[1] ;
 wire \wb_cross_clk.m_wb_i_dat[2] ;
 wire \wb_cross_clk.m_wb_i_dat[3] ;
 wire \wb_cross_clk.m_wb_i_dat[4] ;
 wire \wb_cross_clk.m_wb_i_dat[5] ;
 wire \wb_cross_clk.m_wb_i_dat[6] ;
 wire \wb_cross_clk.m_wb_i_dat[7] ;
 wire \wb_cross_clk.m_wb_i_dat[8] ;
 wire \wb_cross_clk.m_wb_i_dat[9] ;
 wire \wb_cross_clk.msy_xor_ack ;
 wire \wb_cross_clk.msy_xor_err ;
 wire \wb_cross_clk.prev_ack ;
 wire \wb_cross_clk.prev_stb ;
 wire \wb_cross_clk.prev_xor_ack ;
 wire \wb_cross_clk.prev_xor_err ;
 wire \wb_cross_clk.prev_xor_newreq ;
 wire \wb_cross_clk.s_burst_cnt[0] ;
 wire \wb_cross_clk.s_burst_cnt[1] ;
 wire \wb_cross_clk.s_burst_cnt[2] ;
 wire \wb_cross_clk.s_burst_cnt[3] ;
 wire \wb_cross_clk.s_m_sync.d_xfer_xor_sync[0] ;
 wire \wb_cross_clk.s_m_sync.d_xfer_xor_sync[1] ;
 wire \wb_cross_clk.s_m_sync.d_xfer_xor_sync[2] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[0] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[10] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[11] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[12] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[13] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[14] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[15] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[16] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[17] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[1] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[2] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[3] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[4] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[5] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[6] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[7] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[8] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[9] ;
 wire \wb_cross_clk.s_m_sync.s_xfer_xor_flag ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__I (.I(_1522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__I (.I(_1524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__I (.I(_1526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__A1 (.I(_1527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__I (.I(net237),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__A1 (.I(_1527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1608__I (.I(net236),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__A1 (.I(_1527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__I (.I(net235),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1612__A1 (.I(_1527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__I (.I(net234),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A1 (.I(_1527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__I (.I(_1538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__I (.I(_1539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__I (.I(_1526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1621__A1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A1 (.I(_1524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__I (.I(_1543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__I (.I(_1544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1626__A1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__A1 (.I(_1524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1629__I (.I(_1547_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__I (.I(_1548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__A1 (.I(_1527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1634__I (.I(_1551_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1635__I (.I(_1552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1637__I (.I(_1553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__A2 (.I(net25),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__I (.I(_1522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__I1 (.I(net26),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__S (.I(_1557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__A1 (.I(_1526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__C (.I(_1558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__I1 (.I(net8),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__I1 (.I(net9),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__S (.I(_1522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__A1 (.I(_1560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__I1 (.I(net24),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__S (.I(_1557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1647__I1 (.I(net23),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A1 (.I(_1563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A2 (.I(_1564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__I (.I(net90),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__I1 (.I(net7),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__S (.I(_1522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1651__A2 (.I(_1567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__I1 (.I(net6),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__I1 (.I(net17),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__I1 (.I(net16),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A1 (.I(_1570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A2 (.I(_1571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A3 (.I(_1572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1657__I1 (.I(net10),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1657__S (.I(_1557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__I0 (.I(\m_arbiter.wb0_adr[18] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__I1 (.I(net12),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__S (.I(_1557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A1 (.I(_1526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A2 (.I(net18),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__I1 (.I(net15),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1663__A1 (.I(_1526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1663__C (.I(_1579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__I1 (.I(net5),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__S (.I(_1557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__I1 (.I(net4),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__S (.I(_1557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__I1 (.I(net13),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__S (.I(_1557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__I1 (.I(net11),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__S (.I(_1557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__A1 (.I(_1581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__A2 (.I(_1582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__B (.I(net90),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1671__I1 (.I(net14),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__I (.I(_1588_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__I1 (.I(net3),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__A1 (.I(net128),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__A2 (.I(net127),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__I1 (.I(net22),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__S (.I(_1557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__I1 (.I(net21),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__S (.I(_1522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__I (.I(net131),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__A2 (.I(net132),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__A3 (.I(_1593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__I1 (.I(net18),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A1 (.I(_0391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A2 (.I(_1579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1685__A1 (.I(_1571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1685__A2 (.I(_1572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__A1 (.I(_1560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__A3 (.I(_1567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__I1 (.I(net25),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__S (.I(_1557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A1 (.I(_0396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A2 (.I(_1558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A3 (.I(_1581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A4 (.I(_1582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__I1 (.I(net20),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__S (.I(_1522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1691__I (.I(_0398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__I1 (.I(net19),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A1 (.I(net130),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A2 (.I(net129),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A1 (.I(_1570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1696__A2 (.I(_1594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__A1 (.I(_1570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1699__A1 (.I(_1563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1699__A2 (.I(_1564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__I (.I(net132),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__A1 (.I(_0405_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__A3 (.I(_1593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__I (.I(net128),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__A2 (.I(net127),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__A1 (.I(_0403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__A4 (.I(_0409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__I (.I(_0412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__I (.I(_1553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1710__A2 (.I(_0415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__A1 (.I(_1554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__B (.I(_0413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__A1 (.I(_0391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__A2 (.I(_1579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__A1 (.I(_0405_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__A2 (.I(_1570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__A1 (.I(_0391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__A2 (.I(_1579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A1 (.I(\iram_latched[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A2 (.I(_0426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__I (.I(_1553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__A2 (.I(_0415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__A1 (.I(_0428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__B (.I(_0413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__A1 (.I(\iram_latched[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__A2 (.I(_0426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__A2 (.I(_0415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A1 (.I(_0428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A2 (.I(\wb_compressor.wb_i_dat[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__B (.I(_0412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__A1 (.I(\iram_latched[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__A2 (.I(_0426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__A2 (.I(_0436_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__A2 (.I(_0415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__A1 (.I(_0428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__B (.I(_0412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A1 (.I(\iram_latched[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A2 (.I(_0426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__A2 (.I(_0440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A2 (.I(_0415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__A1 (.I(_0428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__A2 (.I(\wb_compressor.wb_i_dat[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__B (.I(_0412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__A1 (.I(\iram_latched[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__A2 (.I(_0426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A2 (.I(_0444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__A2 (.I(_0415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__A1 (.I(_0428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__B (.I(_0412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A1 (.I(\iram_latched[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A2 (.I(_0426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A2 (.I(_0448_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__A2 (.I(_0415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__A1 (.I(_0428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__B (.I(_0412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A1 (.I(\iram_latched[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A2 (.I(_0426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__A2 (.I(_0415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__A1 (.I(_0428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__B (.I(_0412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__A1 (.I(\iram_latched[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__A2 (.I(_0426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1759__I (.I(_0426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1760__I (.I(_1553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__S (.I(_0458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__A1 (.I(\iram_latched[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__A2 (.I(_0457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__B2 (.I(_0413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A2 (.I(_1594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__I (.I(net127),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__A1 (.I(net128),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A1 (.I(net128),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1769__A1 (.I(_1526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A1 (.I(_1524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A2 (.I(net6),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__A1 (.I(net130),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__A2 (.I(net129),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A1 (.I(_0468_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A2 (.I(_0403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__A2 (.I(_0471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__A1 (.I(_0405_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__A3 (.I(net131),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A2 (.I(_0403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A2 (.I(_0403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A4 (.I(_0409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__A2 (.I(net228),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__B1 (.I(net224),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A1 (.I(_0462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A1 (.I(_0460_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A2 (.I(_0478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__S (.I(_0458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A1 (.I(\iram_latched[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A2 (.I(_0457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__B2 (.I(_0413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__A2 (.I(_0471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__A1 (.I(_0462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__A2 (.I(_0483_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__S (.I(_0458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A1 (.I(\iram_latched[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A2 (.I(_0457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__B2 (.I(_0413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A2 (.I(_0471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A1 (.I(_0462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A2 (.I(_0489_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__S (.I(_0458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A1 (.I(\iram_latched[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A2 (.I(_0457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__B2 (.I(_0413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1798__A2 (.I(_0471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__A1 (.I(_0462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__A2 (.I(_0495_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A1 (.I(_0492_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__S (.I(_0458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A2 (.I(_0457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__B2 (.I(_0413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A2 (.I(_0471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__A1 (.I(_0462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__A2 (.I(_0501_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__A1 (.I(_0498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__S (.I(_0458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A2 (.I(_0457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__B2 (.I(_0413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__A2 (.I(_0471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A1 (.I(_0462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A2 (.I(_0507_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A1 (.I(_0504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__S (.I(_0458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A1 (.I(\iram_latched[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A2 (.I(_0457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__B2 (.I(_0413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__A2 (.I(_0471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1822__A1 (.I(_0462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1822__A2 (.I(_0513_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1823__A1 (.I(_0510_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__S (.I(_0415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__A1 (.I(\iram_latched[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__A2 (.I(_0457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__B2 (.I(_0413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__A2 (.I(_0471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__A1 (.I(_0462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__A2 (.I(_0519_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__A1 (.I(_0520_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__A2 (.I(_0516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1831__I (.I(\wb_compressor.wb_ack ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A1 (.I(_1524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A2 (.I(\m_arbiter.i_wb0_cyc ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__A1 (.I(_1526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__A2 (.I(net27),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__B (.I(_0524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__A1 (.I(_1524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__A2 (.I(net46),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A1 (.I(_0525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A2 (.I(_0526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A1 (.I(_1553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A2 (.I(_0527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__B (.I(_0529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A1 (.I(_0521_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A2 (.I(_0412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__A1 (.I(\wb_compressor.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__A1 (.I(net85),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__A2 (.I(net84),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__I (.I(net193),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__I (.I(_0542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__I (.I(_0543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__B (.I(_0544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__A1 (.I(net84),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__B (.I(_0544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__I (.I(_0543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__I (.I(\wb_compressor.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__A1 (.I(_0549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__I (.I(_0542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__I (.I(net84),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__I (.I(_0555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__B (.I(_0556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1871__A1 (.I(_0553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__I (.I(_0558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__S (.I(_0559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__S (.I(_0559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__S (.I(_0559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__A1 (.I(_0560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__S (.I(_0559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__I1 (.I(_1579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__S (.I(_0558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1880__S (.I(_0558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__I1 (.I(_0391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__S (.I(_0559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__A1 (.I(_0564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__A2 (.I(_0565_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__A3 (.I(_0566_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__S (.I(_0558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__S (.I(_0558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__I1 (.I(_1571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__S (.I(_0558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1886__S (.I(_0559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__A1 (.I(_0569_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__A3 (.I(_0571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__A4 (.I(_0572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__A2 (.I(_0575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__A2 (.I(_0542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__I (.I(\sspi.state[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__I (.I(_0524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__I (.I(_0579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__A1 (.I(_0426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__A2 (.I(_0527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__A1 (.I(_1553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__A1 (.I(\wb_compressor.wb_err ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__A2 (.I(_1553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__A1 (.I(_0403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__A4 (.I(_0409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1904__A1 (.I(_0462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__A1 (.I(_0525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__A2 (.I(_0526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__B2 (.I(_0462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A1 (.I(_1553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A1 (.I(\wb_compressor.wb_ack ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A2 (.I(_1553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__S (.I(_0412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__A1 (.I(_0590_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__A2 (.I(_0596_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A1 (.I(_0582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A2 (.I(_0597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__A1 (.I(_0524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__A2 (.I(_0582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1920__A2 (.I(net259),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A1 (.I(_0603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A2 (.I(_0607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__B (.I(\sspi.bit_cnt[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__I (.I(\sspi.bit_cnt[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A1 (.I(_0609_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A2 (.I(_0610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A3 (.I(net259),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1927__A2 (.I(_0611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1929__A2 (.I(_0582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__A1 (.I(_0524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__A2 (.I(_0580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__I (.I(net92),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1936__A1 (.I(_0619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__I (.I(_0524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__I (.I(_0622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__C (.I(_0623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__A1 (.I(_0623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A1 (.I(\sspi.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__I (.I(_0619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A2 (.I(_0629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A3 (.I(_0582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__I (.I(_0579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__B (.I(_0631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A1 (.I(_0622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__A1 (.I(\sspi.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__I (.I(_0579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__A2 (.I(_0611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__A3 (.I(_0636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__A1 (.I(_0582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__B2 (.I(_0639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1961__A1 (.I(_0634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__I (.I(_0622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A1 (.I(_0641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__A1 (.I(_0641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__A2 (.I(_0639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__S (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__I1 (.I(net43),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__S (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__S (.I(_1526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__S (.I(_1526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__I1 (.I(net31),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__S (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__I0 (.I(\m_arbiter.wb0_o_dat[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__S (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__I0 (.I(\m_arbiter.wb0_o_dat[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__S (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__I0 (.I(\m_arbiter.wb0_o_dat[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__S (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A1 (.I(_1526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A2 (.I(net47),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__A1 (.I(_1524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__A2 (.I(_0656_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__A1 (.I(_0457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__A2 (.I(_0658_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__I (.I(_0659_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__I (.I(_0542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A1 (.I(_0660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A3 (.I(_0575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A1 (.I(_0543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__A2 (.I(_0596_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A2 (.I(_0590_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__A1 (.I(_0575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A1 (.I(\wb_compressor.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A3 (.I(_0555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__A1 (.I(\wb_compressor.wb_ack ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__A2 (.I(\wb_compressor.wb_err ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__I (.I(_0676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__A1 (.I(_0521_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A2 (.I(_0677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__A1 (.I(_0677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A1 (.I(\wb_compressor.wb_err ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A2 (.I(_0677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__A1 (.I(_0677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__A2 (.I(net245),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__S (.I(_0677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__S (.I(_0677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__S (.I(_0677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__S (.I(_0677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__S (.I(_0677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__S (.I(_0677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__I (.I(_0676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__S (.I(_0688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2039__S (.I(_0688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__S (.I(_0688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__S (.I(_0688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__S (.I(_0688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__I0 (.I(\wb_compressor.wb_i_dat[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__S (.I(_0688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__S (.I(_0688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__I0 (.I(\wb_compressor.wb_i_dat[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__S (.I(_0688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__S (.I(_0688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__S (.I(_0688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__I (.I(iram_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__A1 (.I(_0700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__A2 (.I(_0457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__A4 (.I(_0596_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__I (.I(_0701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__A1 (.I(_0700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__A2 (.I(\iram_latched[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__I (.I(iram_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A2 (.I(net48),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__B (.I(_0631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2065__A1 (.I(_0700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2065__A2 (.I(\iram_latched[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__A2 (.I(net55),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__B (.I(_0631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__A1 (.I(_0700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__A2 (.I(net56),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__B (.I(_0631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__A1 (.I(_0700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__B (.I(_0631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__A1 (.I(_0700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__A2 (.I(\iram_latched[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__B (.I(_0631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__A1 (.I(_0700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__A2 (.I(\iram_latched[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__B (.I(_0631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__A1 (.I(_0700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__A2 (.I(\iram_latched[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__B (.I(_0631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__A2 (.I(\iram_latched[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__B (.I(_0631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__A2 (.I(\iram_latched[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__I (.I(_0579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__B (.I(_0721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__A2 (.I(\iram_latched[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A1 (.I(iram_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__B (.I(_0721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__A2 (.I(\iram_latched[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__A1 (.I(iram_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__B (.I(_0721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__A2 (.I(\iram_latched[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__A1 (.I(iram_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__B (.I(_0721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A2 (.I(\iram_latched[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__A1 (.I(iram_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__B (.I(_0721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A2 (.I(\iram_latched[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__A1 (.I(iram_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__B (.I(_0721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__A2 (.I(\iram_latched[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__A1 (.I(iram_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2107__B (.I(_0721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__A1 (.I(\iram_latched[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__A2 (.I(_0700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__B (.I(_0721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__A1 (.I(_0700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__A2 (.I(_0631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__S0 (.I(_0737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__S1 (.I(\clk_div.curr_div[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__S0 (.I(_0737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__S1 (.I(\clk_div.curr_div[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__A2 (.I(_0740_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__S0 (.I(_0737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__S1 (.I(\clk_div.curr_div[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2121__S0 (.I(_0737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2121__S1 (.I(\clk_div.curr_div[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__A2 (.I(net244),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__A1 (.I(_1570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__A3 (.I(_0409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A2 (.I(_0525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A3 (.I(_0656_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A2 (.I(_0751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__A1 (.I(_1552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__A2 (.I(_0751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__A2 (.I(_0751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2132__A1 (.I(_1548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2132__A2 (.I(_0751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A2 (.I(_0751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__A1 (.I(_1544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__A2 (.I(_0751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__A2 (.I(_0751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__A1 (.I(_1539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__A2 (.I(_0751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A2 (.I(_0756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__A1 (.I(_0751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__B (.I(_0721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__A1 (.I(_0737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__A2 (.I(_0759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__I (.I(_0622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__A2 (.I(_0759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__C (.I(_0761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__I (.I(\clk_div.curr_div[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2146__I (.I(_0622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__A2 (.I(_0759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__B (.I(_0763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__A2 (.I(_0759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A2 (.I(_0759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__A2 (.I(_0759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__C (.I(_0761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__A2 (.I(_0759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__B (.I(_0763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A2 (.I(_0759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A2 (.I(_0772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__I (.I(_0542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__A2 (.I(_0771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__C (.I(_0774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2162__A2 (.I(_0771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__I (.I(_0776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A2 (.I(_0777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__B (.I(_0544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__A2 (.I(_0776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__A2 (.I(_0777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__C (.I(_0774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A2 (.I(_0771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__A2 (.I(_0777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__B (.I(_0544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__A2 (.I(_0783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A2 (.I(_0777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__B (.I(_0544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__A2 (.I(_0783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__A2 (.I(_0777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__B (.I(_0544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__A2 (.I(_0783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__A2 (.I(_0777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__B (.I(_0544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__A2 (.I(_0783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__A2 (.I(_0777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__B (.I(_0544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__A2 (.I(_0783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A2 (.I(_0777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__I (.I(_0543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__B (.I(_0794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__A1 (.I(\wb_cross_clk.m_s_sync.d_data[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__A2 (.I(_0783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A2 (.I(_0777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__B (.I(_0794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A1 (.I(\wb_cross_clk.m_s_sync.d_data[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A2 (.I(_0783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__A2 (.I(_0777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2195__B (.I(_0794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A1 (.I(\wb_cross_clk.m_s_sync.d_data[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A2 (.I(_0783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__I (.I(_0776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__A2 (.I(_0800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2199__B (.I(_0794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A2 (.I(_0783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__A2 (.I(_0800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__B (.I(_0794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A2 (.I(_0783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__A2 (.I(_0800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2205__B (.I(_0794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A2 (.I(_0806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A2 (.I(_0800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__B (.I(_0794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__A2 (.I(_0806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__A2 (.I(_0800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__B (.I(_0794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__A2 (.I(_0806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A2 (.I(_0800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__B (.I(_0794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__A2 (.I(_0806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A2 (.I(_0800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__B (.I(_0794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__A2 (.I(_0806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__A2 (.I(_0800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__I (.I(_0543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__B (.I(_0817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A2 (.I(_0772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A2 (.I(_0771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__C (.I(_0774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A2 (.I(_0772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__A2 (.I(_0771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__C (.I(_0774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A2 (.I(_0772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A2 (.I(_0771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__C (.I(_0660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A2 (.I(_0806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A2 (.I(_0800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__B (.I(_0817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A2 (.I(_0806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A2 (.I(_0800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__B (.I(_0817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A2 (.I(_0806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__I (.I(_0776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A2 (.I(_0829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__B (.I(_0817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__A2 (.I(_0806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A2 (.I(_0829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__B (.I(_0817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__A2 (.I(_0806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__A2 (.I(_0829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__B (.I(_0817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__A2 (.I(_0835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A2 (.I(_0829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__B (.I(_0817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__A2 (.I(_0835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A2 (.I(_0829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__B (.I(_0817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__A2 (.I(_0835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__A2 (.I(_0829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__B (.I(_0817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__A2 (.I(_0835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__A2 (.I(_0829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__B (.I(_0817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__A2 (.I(_0835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A2 (.I(_0829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__I (.I(_0543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__B (.I(_0846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A2 (.I(_0835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__A2 (.I(_0829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__B (.I(_0846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__A2 (.I(_0835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__A2 (.I(_0829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__B (.I(_0846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A2 (.I(_0835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__I (.I(_0776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__A2 (.I(_0852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__B (.I(_0846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__A2 (.I(_0835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A2 (.I(_0852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__B (.I(_0846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__A2 (.I(_0835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A2 (.I(_0852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__B (.I(_0846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A2 (.I(_0772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A2 (.I(_0852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__B (.I(_0846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A2 (.I(_0852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__A2 (.I(_0771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__B (.I(_0846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2287__A2 (.I(_0776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A2 (.I(_0771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__B (.I(_0846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A2 (.I(_0772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A2 (.I(_0852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__B (.I(_0846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A2 (.I(_0776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__A2 (.I(_0771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__B (.I(_0549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A2 (.I(_0776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A2 (.I(_0771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__B (.I(_0549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A2 (.I(_0772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A2 (.I(_0852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__B (.I(_0549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__A2 (.I(_0772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A2 (.I(_0852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__B (.I(_0549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A2 (.I(_0772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__A2 (.I(_0852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__B (.I(_0549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A2 (.I(_0772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A2 (.I(_0852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__B (.I(_0549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A1 (.I(_0634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A2 (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A2 (.I(\m_arbiter.i_wb0_cyc ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__B (.I(_0412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__C (.I(_0526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__B (.I(_0880_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__C (.I(_0883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__A2 (.I(_0885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A1 (.I(_0634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A2 (.I(_0544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A1 (.I(_0553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A1 (.I(_0553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__I (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A2 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A2 (.I(_0891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__B (.I(_0721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A2 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A2 (.I(_0891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__I (.I(_0579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__B (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__I (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__A2 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__A2 (.I(_0891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__B (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A2 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A2 (.I(_0891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__B (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A2 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A2 (.I(_0891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__B (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A2 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A2 (.I(_0891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__B (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__A2 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A2 (.I(_0891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__B (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__A2 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__A2 (.I(_0891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__B (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A2 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__A2 (.I(_0891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__B (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__A2 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__A2 (.I(_0891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__B (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__A2 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A2 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__C (.I(_0580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__A2 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__A2 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__C (.I(_0580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A2 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A2 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__C (.I(_0580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A2 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__I (.I(_0579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A2 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__C (.I(_0917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A2 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A2 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__C (.I(_0917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__A2 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__A2 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__C (.I(_0917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A2 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A2 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__C (.I(_0917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__A2 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A2 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__C (.I(_0917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__S (.I(_0923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__I (.I(_0885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__A1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A2 (.I(_0925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A1 (.I(_0925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A2 (.I(_0926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A1 (.I(_1527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A2 (.I(net1),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__A2 (.I(_0925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__I1 (.I(_0929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__S (.I(_0923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__I1 (.I(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__S (.I(_0923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__I (.I(_0885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A2 (.I(_0925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A1 (.I(_0933_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A2 (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__A2 (.I(_0925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A1 (.I(_1552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A2 (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__I (.I(_0885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A2 (.I(_0937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A1 (.I(_1548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A2 (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__A2 (.I(_0937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__A1 (.I(_1544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__A2 (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A2 (.I(_0937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__A1 (.I(_1539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__A2 (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A2 (.I(_0937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A1 (.I(net234),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A2 (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__A2 (.I(_0937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A1 (.I(net235),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A2 (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A2 (.I(_0937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__A1 (.I(net236),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__A2 (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A2 (.I(_0937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A1 (.I(net237),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A2 (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__I1 (.I(net148),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__S (.I(_0923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__I1 (.I(net149),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__S (.I(_0923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__I1 (.I(net135),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__S (.I(_0923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__I1 (.I(net136),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__S (.I(_0923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__I1 (.I(net137),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__S (.I(_0949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__I1 (.I(net138),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__S (.I(_0949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__I1 (.I(net139),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__S (.I(_0949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__I1 (.I(net140),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__S (.I(_0949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A2 (.I(_0937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A2 (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A2 (.I(_0937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__A2 (.I(_0925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__I1 (.I(net129),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__S (.I(_0949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__I1 (.I(net130),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__S (.I(_0949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A2 (.I(_0937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A1 (.I(_1593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A2 (.I(_0925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A2 (.I(_0923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__A2 (.I(_0925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__I1 (.I(_1564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__S (.I(_0949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__I1 (.I(_1563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__S (.I(_0949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__I1 (.I(_0396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__S (.I(_0949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__I1 (.I(_1558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__S (.I(_0949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__I1 (.I(_1582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__S (.I(_0964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__I1 (.I(_1581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__S (.I(_0964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A2 (.I(_0923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__A1 (.I(_0468_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__A2 (.I(_0925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__I1 (.I(_1567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__S (.I(_0964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__I1 (.I(_1560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__S (.I(_0964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__S (.I(_0964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__S (.I(_0964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__S (.I(_0964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__S (.I(_0964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__S (.I(_0964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__I1 (.I(_1579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__S (.I(_0964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__I1 (.I(_1572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__S (.I(_0885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__I1 (.I(_1571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__S (.I(_0885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__I1 (.I(_0391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__S (.I(_0885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__I1 (.I(_0525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__S (.I(_0885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A2 (.I(_0676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A1 (.I(_0553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A2 (.I(_0623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A1 (.I(_0623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A2 (.I(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__I (.I(_0982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A1 (.I(_0623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__A1 (.I(_0634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__A2 (.I(_0880_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A2 (.I(_0623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A1 (.I(_0634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__A2 (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A2 (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__B (.I(_0885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__I (.I(_0524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A1 (.I(_1527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A2 (.I(net1),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A1 (.I(_0933_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A1 (.I(_0926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__B (.I(_0988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A3 (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A2 (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__B (.I(_0579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__C (.I(_0925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__A1 (.I(_0933_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__A2 (.I(_0926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A1 (.I(_0923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__A1 (.I(_0623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__A1 (.I(_0926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__B2 (.I(_0885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A1 (.I(_0623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A1 (.I(\wb_compressor.wb_ack ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A2 (.I(\wb_compressor.wb_err ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A1 (.I(_0933_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A1 (.I(_0676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__B (.I(_0549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__B (.I(_0549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A1 (.I(_0543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A1 (.I(\wb_compressor.wb_ack ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A2 (.I(\wb_compressor.wb_err ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__C (.I(_0660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__B (.I(_0676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__A1 (.I(_0553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(_0553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A1 (.I(_0553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__A2 (.I(_0623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A2 (.I(_0544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A1 (.I(\wb_compressor.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A1 (.I(_0542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A2 (.I(_0575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A2 (.I(_0458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A1 (.I(_1554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A2 (.I(_0933_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__A1 (.I(_1027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__A2 (.I(_1029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__A2 (.I(_1027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A2 (.I(_1553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__A1 (.I(_0415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__A2 (.I(_0926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__I (.I(_0559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__A2 (.I(_1033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__A1 (.I(_1033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__A1 (.I(net487),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__A2 (.I(net220),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__B (.I(_1027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A2 (.I(_1027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__I1 (.I(net487),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__S (.I(_1027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A1 (.I(_0542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__I (.I(net213),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__S (.I(_1039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__S (.I(_1039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__I1 (.I(net69),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__S (.I(_1039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__I1 (.I(net70),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__S (.I(_1039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__S (.I(_1039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__S (.I(_1039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__S (.I(_1039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__S (.I(_1039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__S (.I(_1039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__S (.I(_1039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__I1 (.I(net78),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__S (.I(net213),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__I0 (.I(\wb_compressor.wb_i_dat[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__I1 (.I(net79),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__I1 (.I(net80),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__I0 (.I(\wb_compressor.wb_i_dat[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__I1 (.I(net81),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__I1 (.I(net82),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__S (.I(net214),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__I1 (.I(net83),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__S (.I(net214),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__A1 (.I(\wb_compressor.wb_err ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__B2 (.I(net85),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A2 (.I(\wb_compressor.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A3 (.I(_0543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A1 (.I(\wb_compressor.wb_ack ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__B2 (.I(net84),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A2 (.I(\wb_compressor.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A3 (.I(_0543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A1 (.I(_0641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__A1 (.I(_0641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A1 (.I(_0641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A1 (.I(_0634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A2 (.I(\wb_compressor.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__A1 (.I(net250),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A1 (.I(net250),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__B (.I(_0549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__A1 (.I(_0575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__B (.I(net202),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A1 (.I(_0543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A1 (.I(\wb_compressor.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__B1 (.I(_0575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__I (.I(_1554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__I (.I(_0458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A2 (.I(_1074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A1 (.I(_1073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A1 (.I(_0555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A2 (.I(_1077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__I (.I(_1078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__I (.I(_1033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A2 (.I(_1080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__B (.I(_1077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A1 (.I(_1080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A2 (.I(_1552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A1 (.I(_0556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__B (.I(_1079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A1 (.I(net176),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A2 (.I(_1084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__A1 (.I(_1072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__C (.I(_0660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__I (.I(_1077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A1 (.I(net141),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A2 (.I(_1086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__B1 (.I(_1079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__B2 (.I(_0929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A2 (.I(_0458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__A1 (.I(_1554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A2 (.I(_1077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__B1 (.I(_1078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A1 (.I(_0555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__B2 (.I(_1074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__A1 (.I(_1073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__C (.I(_1093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A1 (.I(net177),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A2 (.I(_1072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A1 (.I(_0553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A1 (.I(net142),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A2 (.I(_1086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__B1 (.I(_1079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__B2 (.I(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__I1 (.I(net534),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__S (.I(_0559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__A2 (.I(_1077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__B1 (.I(_1078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__A1 (.I(_0555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__B2 (.I(_1074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__A1 (.I(_1073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__C (.I(_1093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__A1 (.I(net178),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__A2 (.I(_1072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A1 (.I(_0553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__A1 (.I(_1073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__A2 (.I(_1080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__B (.I(_0556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A1 (.I(\wb_cross_clk.m_s_sync.d_data[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A2 (.I(_0428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A1 (.I(_1554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A2 (.I(_1539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A1 (.I(_1029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A2 (.I(_1079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__B2 (.I(_1086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__C (.I(_1093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A1 (.I(net179),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A2 (.I(_1072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__A1 (.I(_0553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A1 (.I(_1033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A2 (.I(_1593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A2 (.I(_1080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__B (.I(_0555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A1 (.I(\wb_cross_clk.m_s_sync.d_data[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A2 (.I(_0428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__A1 (.I(_1074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__A2 (.I(net234),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A1 (.I(net487),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A2 (.I(_1079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__B2 (.I(_1086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A1 (.I(_1093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__A1 (.I(net180),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__A2 (.I(_1084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__A1 (.I(_0774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A1 (.I(_1033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A2 (.I(_1080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__B (.I(_0555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__A1 (.I(\wb_cross_clk.m_s_sync.d_data[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__A2 (.I(_0428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A1 (.I(_1554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A2 (.I(net235),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A1 (.I(net220),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A2 (.I(_1079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__B2 (.I(_1086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A1 (.I(_1093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A1 (.I(net181),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A2 (.I(_1084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__B (.I(_1122_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__A1 (.I(_0774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A2 (.I(_1074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__A1 (.I(_1073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__A2 (.I(net236),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__I1 (.I(net504),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__S (.I(_1033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A1 (.I(_1086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__B2 (.I(_0556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A1 (.I(net182),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A2 (.I(_1084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A1 (.I(_1072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__C (.I(_0660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__A2 (.I(_1074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A1 (.I(_1073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A2 (.I(net237),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__S (.I(_1033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A1 (.I(_1086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__B2 (.I(_0556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A1 (.I(net183),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A2 (.I(_1084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__A1 (.I(_1072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__C (.I(_0660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A1 (.I(_1073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A2 (.I(_1080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__B (.I(_0556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__I1 (.I(net148),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__S (.I(_1033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__A1 (.I(_0564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__A2 (.I(_1078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__B2 (.I(_1086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__C (.I(_1093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A1 (.I(net184),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A2 (.I(_1084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__A1 (.I(_0774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A1 (.I(_1073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A2 (.I(net512),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__A2 (.I(_1080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__B (.I(_0556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__I1 (.I(net149),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__S (.I(_1033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A1 (.I(_0569_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A2 (.I(_1078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__B1 (.I(_1142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__B2 (.I(_1086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2703__C (.I(_1093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__A1 (.I(net185),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__A2 (.I(_1084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A1 (.I(_0774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A1 (.I(_1073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__A2 (.I(_1080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__B (.I(_0555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__I1 (.I(net135),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__S (.I(_0559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A1 (.I(_0566_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A2 (.I(_1078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__B1 (.I(_1148_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__B2 (.I(_1086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__A1 (.I(net187),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__A2 (.I(_1084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__A1 (.I(_0774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__A1 (.I(_1073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__A2 (.I(net515),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__A2 (.I(_1080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__B (.I(_0555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__I1 (.I(net136),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__S (.I(_0559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__A1 (.I(_0560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__A2 (.I(_1078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__B1 (.I(_1154_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__B2 (.I(_1077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__C (.I(_1071_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__A1 (.I(net188),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__A2 (.I(_1084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__A1 (.I(_0774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A2 (.I(\wb_compressor.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__A1 (.I(_1554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__A2 (.I(net137),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__A2 (.I(_1033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__A1 (.I(_1074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__A2 (.I(_1080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__B (.I(_0555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A1 (.I(_1158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A3 (.I(_1160_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A1 (.I(_0565_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A2 (.I(_1079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__A1 (.I(net189),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__A2 (.I(_1084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__A1 (.I(_1072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__C (.I(_0660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A1 (.I(_1554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A2 (.I(net138),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__A2 (.I(_1074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__B (.I(_1158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A1 (.I(_0556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__B1 (.I(_0572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__B2 (.I(_1079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A1 (.I(net190),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A2 (.I(_1093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__A1 (.I(_1072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__C (.I(_0660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__A1 (.I(_1554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__A2 (.I(net139),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A2 (.I(_1074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__B (.I(_1158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A1 (.I(_0556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__B1 (.I(_0571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__B2 (.I(_1079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__C (.I(_1171_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__A1 (.I(net191),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__A2 (.I(_1093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__A1 (.I(_1072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__C (.I(_0660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__A1 (.I(_1554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__A2 (.I(net140),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__A2 (.I(_1074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__B (.I(_1158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__A1 (.I(_0556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__B2 (.I(_1079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__A1 (.I(net192),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__A2 (.I(_1093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__A1 (.I(_1072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__C (.I(_0660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A1 (.I(\sspi.state[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__A1 (.I(\sspi.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__A1 (.I(_0597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__A1 (.I(_1527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__A2 (.I(_0590_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__C (.I(_0917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__A1 (.I(\sspi.state[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__A1 (.I(\sspi.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__A2 (.I(_0639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__A1 (.I(\sspi.state[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__A2 (.I(\sspi.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A1 (.I(_0639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__A1 (.I(_0597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__B (.I(_0641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A1 (.I(_1200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A2 (.I(_0607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__B (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__A1 (.I(_1202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__B (.I(_0603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__B (.I(_1202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__A1 (.I(_0603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__I (.I(_0579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__B (.I(_1207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__I (.I(\sspi.bit_cnt[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__A1 (.I(_0610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__A2 (.I(net259),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__A1 (.I(_1200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__A1 (.I(_1208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__A1 (.I(_0609_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__B2 (.I(_0639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2783__A1 (.I(_1208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A1 (.I(_0634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A1 (.I(_0639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A2 (.I(_0636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__A1 (.I(\sspi.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__A1 (.I(_0639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__B (.I(_1207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__A3 (.I(_0639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__A1 (.I(_0582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__A2 (.I(_0597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__I (.I(_1223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__A2 (.I(_1224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A1 (.I(_0516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A2 (.I(_0520_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A3 (.I(_1223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A1 (.I(_0988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__I (.I(_1223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A1 (.I(_0510_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A3 (.I(_1227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__I (.I(_1223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A2 (.I(_1229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__B (.I(_0641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A1 (.I(_0504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A3 (.I(_1227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A2 (.I(_1229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__B (.I(_0641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__A1 (.I(_0498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__A3 (.I(_1227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__A2 (.I(_1224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__B (.I(_0641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__A1 (.I(_0492_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__A3 (.I(_1227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__A1 (.I(\sspi.res_data[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__A2 (.I(_1224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__B (.I(_0763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2814__A3 (.I(_1227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__A1 (.I(\sspi.res_data[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__A2 (.I(_1224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__B (.I(_0763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__A3 (.I(_1227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A1 (.I(\sspi.res_data[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A2 (.I(_1224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__B (.I(_0763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A1 (.I(_0460_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A2 (.I(_0478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A3 (.I(_1223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__A2 (.I(_1224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__B (.I(_0763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__I (.I(net125),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__A2 (.I(_1224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__A2 (.I(_1229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__C (.I(_0917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2826__I (.I(net126),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2827__A2 (.I(_1224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__A2 (.I(_1229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__C (.I(_0917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2830__A2 (.I(_1224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__A2 (.I(_1229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__C (.I(_0917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A2 (.I(_1224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__A2 (.I(_1229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__C (.I(_0917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__A2 (.I(_1227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__I (.I(_0579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__A2 (.I(_1229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__C (.I(_1253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__A2 (.I(_1227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__A2 (.I(_1229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__C (.I(_1253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__A2 (.I(_1227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__A2 (.I(_1229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__C (.I(_1253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__I (.I(net117),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__A2 (.I(_1227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__A2 (.I(_1229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__C (.I(_1253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__I (.I(net92),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A1 (.I(\sspi.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A2 (.I(_0582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A1 (.I(_0611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A2 (.I(_1261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__B (.I(_0763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__A1 (.I(_1260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__A2 (.I(_1261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__A2 (.I(_1265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__A1 (.I(_0629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__A3 (.I(net253),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__A2 (.I(net253),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__B (.I(_1207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__A2 (.I(_1270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__A1 (.I(_0629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__A2 (.I(_0611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__A4 (.I(_1271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__A2 (.I(_1271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__B (.I(_1207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A1 (.I(_1200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A1 (.I(_0629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A3 (.I(_1275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A2 (.I(_1275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__B (.I(_1207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__A1 (.I(_1202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__A2 (.I(_0619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__A1 (.I(_1202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__B (.I(_1207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A1 (.I(_1261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__B (.I(_0763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A1 (.I(_1260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A1 (.I(net92),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A2 (.I(_0611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A1 (.I(_1261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__B (.I(_0763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A2 (.I(_0636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A3 (.I(_1261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__B (.I(_0622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A1 (.I(_1260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__A1 (.I(\sspi.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__A2 (.I(_0582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__I (.I(_1294_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__A1 (.I(_0609_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__A2 (.I(_1202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__A3 (.I(_0607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A1 (.I(_1295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__A1 (.I(\sspi.bit_cnt[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__A2 (.I(_0610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__A3 (.I(net259),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A1 (.I(_0619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A2 (.I(_1261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A1 (.I(_0988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A1 (.I(_0619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A2 (.I(_0636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A3 (.I(_1295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__A1 (.I(_1208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__A1 (.I(_1261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__B (.I(\sspi.req_data[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__B (.I(_1207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__A3 (.I(_1270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A1 (.I(_1208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A2 (.I(_1295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A3 (.I(_1271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__A1 (.I(_1295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__A1 (.I(_0634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A1 (.I(_0619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A2 (.I(_0636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A3 (.I(_1275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A1 (.I(_1208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A2 (.I(_1294_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A3 (.I(_1275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__A1 (.I(_1295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__A1 (.I(_0634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__A1 (.I(_0609_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__A2 (.I(_0610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__A3 (.I(_1260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__A4 (.I(_0607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__A1 (.I(_1208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__A2 (.I(_1202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__A3 (.I(net259),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__A4 (.I(_1294_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__A1 (.I(_1295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__A1 (.I(_0634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__A2 (.I(_0636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__A1 (.I(_1260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__A1 (.I(_1295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__A1 (.I(_1261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__B (.I(_1207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2918__A2 (.I(_0636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A1 (.I(_1295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__A1 (.I(_1261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__B (.I(_1207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__A1 (.I(_0629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__A3 (.I(_1295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__A2 (.I(_1295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__B (.I(_1207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__A1 (.I(_0639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__A2 (.I(_0611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__A1 (.I(\sspi.req_addr[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__B (.I(_0622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A1 (.I(_1260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__A1 (.I(_0639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__A2 (.I(net253),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__A2 (.I(_0611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__A2 (.I(_0611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__B (.I(net92),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__A1 (.I(_1208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__A3 (.I(_1265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__A4 (.I(_1332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__A1 (.I(_1331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2940__I (.I(_0579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__B (.I(_1335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__A1 (.I(\sspi.bit_cnt[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__A3 (.I(_1270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__A1 (.I(_1336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__A1 (.I(_0629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__A2 (.I(_1331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__B (.I(_1335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__A1 (.I(\sspi.bit_cnt[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__A2 (.I(_1200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__A1 (.I(_1336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__A1 (.I(_1336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__A2 (.I(_1332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__A1 (.I(_0988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__A1 (.I(\sspi.bit_cnt[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__A2 (.I(_0610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__A3 (.I(_0607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__I0 (.I(_0619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__A1 (.I(_0641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__A2 (.I(_1332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__A1 (.I(_1331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__A2 (.I(_0611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__B (.I(\sspi.req_addr[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__B (.I(_1335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A2 (.I(_0636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A3 (.I(_1270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__A1 (.I(_0629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__A3 (.I(_1331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__B (.I(_1335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A2 (.I(_0636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A3 (.I(_1332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__A3 (.I(_1336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__A1 (.I(_1331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__B2 (.I(\sspi.req_addr[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__A1 (.I(_0580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__A2 (.I(_1336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__B (.I(\sspi.req_addr[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2972__A1 (.I(_0619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__A1 (.I(_0988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__A1 (.I(_0619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__A2 (.I(_0636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__A4 (.I(_1336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__B (.I(_1335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__A1 (.I(_1208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__A2 (.I(_1271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__A3 (.I(_1336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__A2 (.I(_1331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2979__A1 (.I(_0580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__A1 (.I(_1208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__A2 (.I(_1275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__A3 (.I(_1336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A2 (.I(_1331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__A1 (.I(_0580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__A1 (.I(_1208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__A2 (.I(_1202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__A3 (.I(net259),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__A4 (.I(_1336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2984__A2 (.I(_1331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2985__A1 (.I(_0580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__A2 (.I(_1331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__B (.I(\sspi.req_addr[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__B (.I(_1335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__A2 (.I(_1331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2990__B (.I(\sspi.req_addr[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__B (.I(_1335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__A1 (.I(_0629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__A3 (.I(_1336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2993__B (.I(\sspi.req_addr[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__B (.I(_1335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2995__A1 (.I(_0611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__I (.I(_1332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2998__B2 (.I(\sspi.req_addr[16] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__A1 (.I(_0580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3000__B (.I(\sspi.req_addr[17] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3002__A2 (.I(_1380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__B (.I(_1335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__A2 (.I(_1380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A1 (.I(_0629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__B (.I(_0622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__A2 (.I(_1380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__A1 (.I(_1332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__A3 (.I(_1380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__A1 (.I(_0988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__A2 (.I(_1380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__A1 (.I(_0629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__B (.I(_0622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3015__A2 (.I(_1380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__B (.I(_1335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__A2 (.I(_1380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__A1 (.I(_0619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__A1 (.I(_0988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__A2 (.I(_1380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__B2 (.I(\sspi.req_addr[23] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__A1 (.I(_0580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3026__A1 (.I(_0524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__I (.I(_1399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__A1 (.I(\sspi.state[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__A2 (.I(_1399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__I (.I(_1401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__A2 (.I(_1400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__B (.I(_1402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__S (.I(_1402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__S (.I(_1402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__S (.I(_1402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__S (.I(_1402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__S (.I(_1402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__S (.I(_1402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__S (.I(_1402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__S (.I(_1402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__S (.I(_1402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__I0 (.I(\sspi.req_data[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__S (.I(_1401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__S (.I(_1401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__S (.I(_1401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__S (.I(_1401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__I1 (.I(\m_arbiter.wb0_o_dat[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__S (.I(_1401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__I1 (.I(\m_arbiter.wb0_o_dat[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__S (.I(_1401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__I1 (.I(\m_arbiter.wb0_o_dat[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__S (.I(_1401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__I (.I(net244),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__A2 (.I(_1419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__A1 (.I(_1419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__A1 (.I(_1419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3073__A1 (.I(_1419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A1 (.I(_0756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3079__A1 (.I(_1419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__A1 (.I(_1419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__A1 (.I(_1419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__A1 (.I(_1419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3094__A1 (.I(net244),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__B (.I(_0756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__B (.I(_0756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__B (.I(_0756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__B (.I(_0756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3108__A1 (.I(_1419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__A1 (.I(_1419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__A1 (.I(\m_arbiter.i_wb0_cyc ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__B (.I(_0763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3117__A1 (.I(_0597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__A2 (.I(_1200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__B1 (.I(_1265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A2 (.I(_0607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__B1 (.I(_1270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__A1 (.I(_1202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__A1 (.I(\sspi.res_data[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__A2 (.I(net259),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__B2 (.I(\sspi.res_data[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__A2 (.I(_0603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__B2 (.I(\sspi.res_data[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__B (.I(_0610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__A2 (.I(_0603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__A2 (.I(net259),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__B (.I(_1202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__A2 (.I(_1270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__B (.I(_1202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__A2 (.I(_1200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__B1 (.I(_0607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__C1 (.I(_1265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__B (.I(\sspi.bit_cnt[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3130__A1 (.I(\sspi.bit_cnt[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3133__A1 (.I(\sspi.state[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3134__A1 (.I(net195),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A1 (.I(_0761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3136__I1 (.I(\sspi.req_addr[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3136__S (.I(_1400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3138__S (.I(_1400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__S (.I(_1400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3142__S (.I(_1400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__S (.I(_1400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__I (.I(_1399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__I1 (.I(\sspi.req_addr[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__S (.I(_1478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__S (.I(_1478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__I1 (.I(\sspi.req_addr[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__S (.I(_1478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__A1 (.I(\sspi.req_addr[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__A2 (.I(_1400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3154__A2 (.I(_1400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__S (.I(_1478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__S (.I(_1478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__S (.I(_1478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__S (.I(_1478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__I1 (.I(\sspi.req_addr[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__S (.I(_1478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__I1 (.I(\sspi.req_addr[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__S (.I(_1478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__I1 (.I(\sspi.req_addr[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__S (.I(_1478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__I1 (.I(\sspi.req_addr[16] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__S (.I(_1399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__I1 (.I(\sspi.req_addr[17] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__S (.I(_1399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__I0 (.I(\m_arbiter.wb0_adr[18] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__S (.I(_1399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__S (.I(_1399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__S (.I(_1399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__S (.I(_1399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__S (.I(_1399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__A1 (.I(\sspi.req_addr[23] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__A2 (.I(_1400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__A2 (.I(_1400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__A4 (.I(_0658_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__I (.I(_1498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__A2 (.I(_1499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__A1 (.I(_1552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__A2 (.I(_1499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__C (.I(_0761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A2 (.I(_1499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__A1 (.I(_1548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__A2 (.I(_1499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__C (.I(_0761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A2 (.I(_1498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__A1 (.I(_1544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__A2 (.I(_1499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__C (.I(_0761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__A2 (.I(_1498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__A1 (.I(_1539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__A2 (.I(_1499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__C (.I(_0761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__A2 (.I(_1498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__A1 (.I(net234),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__A2 (.I(_1499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__C (.I(_0761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__A2 (.I(_1498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__A1 (.I(net235),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__A2 (.I(_1499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__C (.I(_0761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__A2 (.I(_1498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__A1 (.I(net236),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__A2 (.I(_1499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__C (.I(_0761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__A2 (.I(_1498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__A1 (.I(net237),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__A2 (.I(_1499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__C (.I(_0623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__A3 (.I(net233),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__A4 (.I(_0658_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__I (.I(_1508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__A2 (.I(_1509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__A1 (.I(_1552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__A2 (.I(_1509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__C (.I(_1253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__A2 (.I(_1509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__A1 (.I(_1548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__A2 (.I(_1509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__C (.I(_1253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__A2 (.I(_1508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__A1 (.I(_1544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__A2 (.I(_1509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__C (.I(_1253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__A2 (.I(_1508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__A1 (.I(_1539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__A2 (.I(_1509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__C (.I(_1253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__A2 (.I(_1508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__A1 (.I(net234),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__A2 (.I(_1509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__C (.I(_1253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__A2 (.I(_1508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__A1 (.I(net235),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__A2 (.I(_1509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__C (.I(_1253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__A2 (.I(_1508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__A1 (.I(net236),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__A2 (.I(_1509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__C (.I(_0988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__A2 (.I(_1508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A1 (.I(net237),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A2 (.I(_1509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__C (.I(_0988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__A1 (.I(_1527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__A2 (.I(net27),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__A1 (.I(\m_arbiter.i_wb0_cyc ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__C (.I(_0988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__CLK (.I(clknet_4_2_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__CLK (.I(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__CLK (.I(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__D (.I(net90),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__D (.I(net87),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3245__CLK (.I(clknet_4_14_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__CLK (.I(clknet_4_12_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__CLK (.I(clknet_4_14_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__CLK (.I(clknet_4_15_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__CLK (.I(clknet_4_15_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3250__CLK (.I(clknet_4_11_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__CLK (.I(clknet_4_15_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3252__CLK (.I(clknet_4_15_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__CLK (.I(clknet_4_13_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__CLK (.I(clknet_4_13_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3255__CLK (.I(clknet_4_15_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__CLK (.I(clknet_4_13_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__CLK (.I(clknet_4_5_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__CLK (.I(clknet_4_7_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3259__CLK (.I(clknet_4_5_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__CLK (.I(clknet_4_4_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3261__CLK (.I(clknet_4_7_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__CLK (.I(clknet_4_13_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3263__CLK (.I(clknet_leaf_31_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3268__CLK (.I(clknet_leaf_31_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__CLK (.I(clknet_leaf_31_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3270__CLK (.I(clknet_leaf_31_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__CLK (.I(clknet_4_1_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__CLK (.I(clknet_4_1_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__CLK (.I(clknet_4_1_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3295__CLK (.I(clknet_4_3_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__CLK (.I(clknet_4_8_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__CLK (.I(clknet_4_8_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__CLK (.I(clknet_4_10_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__CLK (.I(clknet_4_10_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__CLK (.I(clknet_4_10_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__CLK (.I(clknet_4_10_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__CLK (.I(clknet_4_10_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__CLK (.I(clknet_4_10_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__CLK (.I(clknet_4_10_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__CLK (.I(clknet_4_11_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3306__CLK (.I(clknet_4_11_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__CLK (.I(clknet_4_11_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__CLK (.I(clknet_4_11_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__CLK (.I(clknet_4_11_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3310__CLK (.I(clknet_4_11_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__CLK (.I(clknet_4_14_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3312__CLK (.I(clknet_4_14_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__CLK (.I(clknet_4_12_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3314__CLK (.I(clknet_4_11_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3315__CLK (.I(clknet_4_8_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__CLK (.I(clknet_4_10_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__CLK (.I(clknet_4_10_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__CLK (.I(clknet_4_10_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__CLK (.I(clknet_4_8_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__CLK (.I(clknet_4_11_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__CLK (.I(clknet_4_8_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__CLK (.I(clknet_4_8_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__CLK (.I(clknet_4_8_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__CLK (.I(clknet_4_6_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__CLK (.I(clknet_4_6_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3328__CLK (.I(clknet_4_6_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__CLK (.I(clknet_4_7_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__CLK (.I(clknet_4_7_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3331__CLK (.I(clknet_4_6_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__CLK (.I(clknet_4_6_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__CLK (.I(clknet_4_6_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__CLK (.I(clknet_4_4_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__CLK (.I(clknet_4_4_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3336__CLK (.I(clknet_4_1_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__CLK (.I(clknet_4_4_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__CLK (.I(clknet_4_1_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__CLK (.I(clknet_leaf_5_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__CLK (.I(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__CLK (.I(clknet_4_3_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__D (.I(_0122_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3343__CLK (.I(clknet_4_8_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__CLK (.I(clknet_leaf_38_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3376__CLK (.I(clknet_leaf_31_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3377__CLK (.I(clknet_leaf_31_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__CLK (.I(clknet_leaf_31_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3381__CLK (.I(clknet_leaf_31_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__CLK (.I(clknet_leaf_31_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__CLK (.I(clknet_leaf_31_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__CLK (.I(clknet_leaf_38_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__CLK (.I(clknet_leaf_38_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3392__CLK (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__CLK (.I(clknet_2_0__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__CLK (.I(clknet_leaf_5_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__CLK (.I(clknet_leaf_5_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__CLK (.I(clknet_leaf_5_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__CLK (.I(clknet_4_1_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__CLK (.I(clknet_leaf_5_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__CLK (.I(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__CLK (.I(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__CLK (.I(clknet_4_1_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__CLK (.I(clknet_4_3_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__CLK (.I(clknet_4_1_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3425__CLK (.I(clknet_4_3_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__CLK (.I(clknet_4_14_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__CLK (.I(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__CLK (.I(clknet_4_2_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__CLK (.I(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__CLK (.I(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__CLK (.I(clknet_4_15_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__CLK (.I(clknet_4_15_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__CLK (.I(clknet_4_15_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__CLK (.I(clknet_4_14_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__CLK (.I(clknet_4_15_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__CLK (.I(clknet_4_15_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__CLK (.I(clknet_4_15_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__CLK (.I(clknet_4_13_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__CLK (.I(clknet_4_13_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__CLK (.I(clknet_4_13_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__CLK (.I(clknet_4_5_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__CLK (.I(clknet_4_5_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__CLK (.I(clknet_4_5_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__CLK (.I(clknet_4_5_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__CLK (.I(clknet_4_7_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__CLK (.I(clknet_4_12_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__CLK (.I(clknet_4_6_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__CLK (.I(clknet_4_6_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__CLK (.I(clknet_4_3_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__CLK (.I(clknet_4_3_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__CLK (.I(clknet_4_14_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__CLK (.I(clknet_4_14_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__CLK (.I(clknet_4_14_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__CLK (.I(clknet_4_12_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__CLK (.I(clknet_4_14_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__CLK (.I(clknet_4_14_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__CLK (.I(clknet_4_12_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__CLK (.I(clknet_4_12_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__CLK (.I(clknet_4_12_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__CLK (.I(clknet_4_12_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__CLK (.I(clknet_4_12_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__CLK (.I(clknet_4_12_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__CLK (.I(clknet_4_2_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__CLK (.I(clknet_4_2_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__CLK (.I(clknet_4_3_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__CLK (.I(clknet_4_3_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__CLK (.I(clknet_4_2_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__CLK (.I(clknet_4_2_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__CLK (.I(clknet_4_3_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__CLK (.I(clknet_leaf_5_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__CLK (.I(clknet_leaf_5_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__CLK (.I(clknet_leaf_16_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__CLK (.I(clknet_leaf_16_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__CLK (.I(clknet_leaf_16_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__CLK (.I(clknet_leaf_16_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__CLK (.I(clknet_leaf_16_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__CLK (.I(clknet_leaf_16_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__CLK (.I(clknet_leaf_8_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__CLK (.I(clknet_leaf_16_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__CLK (.I(clknet_leaf_16_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__CLK (.I(clknet_leaf_9_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__CLK (.I(clknet_leaf_9_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__CLK (.I(clknet_leaf_9_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__CLK (.I(clknet_leaf_8_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__CLK (.I(clknet_leaf_9_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__CLK (.I(clknet_leaf_8_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__CLK (.I(clknet_leaf_8_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__CLK (.I(clknet_leaf_8_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__CLK (.I(clknet_leaf_8_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__CLK (.I(clknet_leaf_9_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__CLK (.I(clknet_leaf_9_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__CLK (.I(clknet_leaf_8_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__CLK (.I(clknet_leaf_8_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__CLK (.I(clknet_leaf_9_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__CLK (.I(clknet_leaf_16_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__CLK (.I(clknet_leaf_5_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__CLK (.I(clknet_leaf_9_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3587__CLK (.I(clknet_leaf_8_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__CLK (.I(clknet_leaf_5_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__CLK (.I(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__CLK (.I(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__CLK (.I(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__CLK (.I(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__I (.I(net249),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__I (.I(net249),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__I (.I(net249),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__I (.I(net249),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__I (.I(net249),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__I (.I(net249),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__I (.I(net249),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__I (.I(net249),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__I (.I(net249),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__I (.I(net249),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__I (.I(net250),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__I (.I(net250),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__I (.I(net250),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__I (.I(net250),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__I (.I(net250),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__I (.I(net250),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_net196_I (.I(net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_user_clock2_I (.I(user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_user_clock2_I (.I(clknet_0_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_user_clock2_I (.I(clknet_0_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_user_clock2_I (.I(clknet_0_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_user_clock2_I (.I(clknet_0_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9_0_net196_I (.I(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_user_clock2_I (.I(clknet_2_0__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_user_clock2_I (.I(clknet_2_0__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_user_clock2_I (.I(clknet_2_3__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_user_clock2_I (.I(clknet_2_3__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_user_clock2_I (.I(clknet_2_3__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_user_clock2_I (.I(clknet_2_3__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_user_clock2_I (.I(clknet_2_3__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_user_clock2_I (.I(clknet_2_3__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_user_clock2_I (.I(clknet_2_3__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_user_clock2_I (.I(clknet_2_3__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_user_clock2_I (.I(clknet_2_3__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_user_clock2_I (.I(clknet_2_0__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_user_clock2_I (.I(clknet_2_3__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_user_clock2_I (.I(clknet_2_3__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_user_clock2_I (.I(clknet_2_3__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_user_clock2_I (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_user_clock2_I (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_user_clock2_I (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_user_clock2_I (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_user_clock2_I (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_user_clock2_I (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_user_clock2_I (.I(clknet_2_0__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_user_clock2_I (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_user_clock2_I (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_user_clock2_I (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_user_clock2_I (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_user_clock2_I (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_user_clock2_I (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_user_clock2_I (.I(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_user_clock2_I (.I(clknet_2_0__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_user_clock2_I (.I(clknet_2_0__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_user_clock2_I (.I(clknet_2_0__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_user_clock2_I (.I(clknet_2_0__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_user_clock2_I (.I(clknet_2_0__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_user_clock2_I (.I(clknet_2_0__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_user_clock2_I (.I(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout249_I (.I(net250),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold106_I (.I(_1563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold109_I (.I(_1570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold114_I (.I(_0396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold117_I (.I(_1564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold120_I (.I(_1567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold122_I (.I(_1582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold125_I (.I(_1558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold128_I (.I(_1581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold131_I (.I(_1560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold134_I (.I(_1572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold141_I (.I(net130),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold147_I (.I(net129),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold99_I (.I(inner_wb_8_burst),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(inner_wb_adr[16]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(inner_wb_adr[17]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(inner_wb_adr[18]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(inner_wb_adr[19]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(inner_wb_adr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(inner_wb_adr[20]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(inner_wb_adr[21]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(inner_wb_adr[22]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(inner_wb_adr[23]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(inner_wb_adr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(inner_wb_4_burst),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(inner_wb_adr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(inner_wb_adr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(inner_wb_adr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(inner_wb_adr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(inner_wb_adr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(inner_wb_adr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(inner_wb_adr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(inner_wb_cyc),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(inner_wb_o_dat[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(inner_wb_o_dat[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(inner_wb_o_dat[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(inner_wb_o_dat[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(inner_wb_o_dat[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(inner_wb_o_dat[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(inner_wb_o_dat[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(inner_wb_o_dat[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(inner_wb_o_dat[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(inner_wb_o_dat[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(inner_wb_o_dat[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(inner_wb_o_dat[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(inner_wb_adr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(inner_wb_o_dat[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(inner_wb_o_dat[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(inner_wb_o_dat[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(inner_wb_o_dat[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(inner_wb_sel[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(inner_wb_sel[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(inner_wb_stb),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(inner_wb_we),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(iram_o_data[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(iram_o_data[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(inner_wb_adr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(iram_o_data[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(iram_o_data[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(iram_o_data[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(iram_o_data[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(iram_o_data[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(iram_o_data[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(iram_o_data[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(iram_o_data[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(iram_o_data[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(iram_o_data[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(inner_wb_adr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(iram_o_data[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(iram_o_data[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(iram_o_data[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(iram_o_data[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(la_data_in[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(la_oenb[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(m_io_in[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(m_io_in[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(m_io_in[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(m_io_in[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(inner_wb_adr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(m_io_in[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(m_io_in[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(m_io_in[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(m_io_in[16]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(m_io_in[17]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(m_io_in[18]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(m_io_in[19]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(m_io_in[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(m_io_in[20]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(m_io_in[21]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(inner_wb_adr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(m_io_in[22]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(m_io_in[23]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(m_io_in[24]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(m_io_in[25]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(m_io_in[26]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(m_io_in[27]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(m_io_in[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(m_io_in[30]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(m_io_in[31]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(m_io_in[32]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(inner_wb_adr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(m_io_in[33]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(m_io_in[34]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(m_io_in[35]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(m_io_in[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(m_io_in[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input95_I (.I(m_io_in[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(m_io_in[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input97_I (.I(m_io_in[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input98_I (.I(mgt_wb_rst_i),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(inner_wb_adr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap208_I (.I(_1071_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap212_I (.I(net213),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap213_I (.I(net214),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap223_I (.I(net224),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap227_I (.I(net228),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap232_I (.I(net233),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output108_I (.I(net392),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output118_I (.I(net118),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net121),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output122_I (.I(net122),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output125_I (.I(net125),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output126_I (.I(net126),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output127_I (.I(net127),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output128_I (.I(net128),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output129_I (.I(net129),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output130_I (.I(net130),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output131_I (.I(net131),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output132_I (.I(net132),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output135_I (.I(net135),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output136_I (.I(net136),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output137_I (.I(net137),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output138_I (.I(net138),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output139_I (.I(net139),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output140_I (.I(net140),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output141_I (.I(net141),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output142_I (.I(net142),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output149_I (.I(net149),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output168_I (.I(net250),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output176_I (.I(net176),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output177_I (.I(net177),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output178_I (.I(net178),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output179_I (.I(net179),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output180_I (.I(net180),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output181_I (.I(net181),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output182_I (.I(net182),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output183_I (.I(net183),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output184_I (.I(net184),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output185_I (.I(net185),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net187),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output188_I (.I(net188),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output189_I (.I(net189),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output190_I (.I(net190),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output191_I (.I(net191),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output192_I (.I(net192),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output193_I (.I(net193),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output195_I (.I(net195),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output196_I (.I(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output202_I (.I(net202),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer1_I (.I(_1522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer2_I (.I(_1522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1_I (.I(net495),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire210_I (.I(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire211_I (.I(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire228_I (.I(_0474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire231_I (.I(net233),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire234_I (.I(_1535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire235_I (.I(_1533_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire236_I (.I(_1531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire237_I (.I(_1529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire241_I (.I(_1594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire260_I (.I(net261),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_145 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_425 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_491 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_509 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_701 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_744 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_490 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_495 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_742 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_829 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_56 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_64 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_421 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_65 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_724 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_75 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_4 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_97 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_357 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_43 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_23 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_25 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_63 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_735 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_806 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_810 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_86 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_25 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_33 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_509 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_794 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_843 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_388 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_4 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_526 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_90 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_145 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_443 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_52 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_705 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_74 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_742 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_83 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_87 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_62 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_670 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_47 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_51 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_62 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_687 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_703 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_39 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_48 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_490 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_565 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_63 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_35 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_99 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_420 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_4 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_40 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_44 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_48 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_530 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_77 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_79 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_145 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_44 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_65 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_724 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_75 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_86 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_38 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_40 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_724 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_736 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_740 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_806 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_821 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_89 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_31 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_56 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_703 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_46 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_742 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_703 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_794 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_703 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_87 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_91 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_687 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_735 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_90 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_4 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_63 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_71 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_724 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_54 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_64 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_392 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_86 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_36 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_40 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_598 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_735 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_794 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_829 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_4 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_495 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_79 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_83 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_99 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_24 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_33 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_38 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_54 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_735 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_829 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_46 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_490 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_54 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_794 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_46 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_62 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_829 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_90 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_408 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_583 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_587 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_674 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_24 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_51 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_670 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_736 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_821 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_828 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_90 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_355 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_408 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_666 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_806 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_828 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_23 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_27 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_79 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_81 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_4 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_44 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_23 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_39 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_443 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_89 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_93 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_97 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_509 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_687 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_87 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_91 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_97 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_36 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_39 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_4 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_526 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_89 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_65 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_75 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_78 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_408 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_52 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_668 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_93 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_24 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_51 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_843 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_845 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_24 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_47 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_526 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_534 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_74 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_90 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_355 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_44 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_392 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_43 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_483 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_99 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_46 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_491 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_54 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_38 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_530 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_534 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_736 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_808 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_89 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_97 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_821 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_38 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_392 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_40 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_47 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_63 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_687 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_806 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_44 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_52 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_56 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_63 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_740 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_392 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_54 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_62 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_86 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_90 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_93 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_97 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_38 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_674 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_808 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_810 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_97 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_39 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_509 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_54 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_724 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_52 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_56 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_74 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_77 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_97 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_4 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_565 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_77 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_79 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_19 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_27 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_31 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_33 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_64 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_740 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_744 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_794 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_808 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_93 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_794 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_93 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_357 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_666 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_814 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_583 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_75 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_829 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_853 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_68 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_78 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_79 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_80 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_81 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_82 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_83 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_84 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_85 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_86 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_87 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_69 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_88 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_89 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_90 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_91 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_92 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_93 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_94 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_95 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_96 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_97 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_98 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_99 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_100 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_102 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_103 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_104 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_106 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_107 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_71 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_109 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_110 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_111 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_112 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_113 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_114 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_115 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_116 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_117 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_72 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_118 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_119 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_120 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_121 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_122 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_123 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_124 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_125 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_126 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_127 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_128 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_129 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_130 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_131 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_132 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_133 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_134 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_135 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_74 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_75 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_76 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_77 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_136 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_138 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_139 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_140 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_142 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_143 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_145 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_146 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_147 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_148 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_149 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_150 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_151 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_152 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_153 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_154 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_155 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_156 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_157 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_158 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_159 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_160 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_269 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_270 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_271 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_272 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_273 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_274 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_275 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_276 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_277 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_278 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_280 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_281 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_282 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_284 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_285 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_287 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_288 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_289 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_290 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_291 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_292 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_293 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_294 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_295 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_296 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_297 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_298 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_299 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_300 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_301 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_302 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_303 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_304 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_305 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_306 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_307 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_308 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_309 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_310 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_311 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_312 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_313 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_315 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_316 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_317 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_319 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_320 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_322 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_323 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_324 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_325 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_326 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_327 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_328 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_329 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_330 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_331 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_332 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_333 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_334 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_335 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_336 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_337 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_338 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_339 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_340 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_341 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_342 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_343 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_344 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_345 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_346 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_347 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_348 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_349 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_351 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_352 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_353 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_355 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_356 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_358 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_359 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_360 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_361 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_362 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_363 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_364 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_365 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_366 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_367 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_368 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_369 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_370 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_371 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_372 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_373 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_374 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_375 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_376 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_377 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_378 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_379 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_380 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_381 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_382 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_383 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_384 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_386 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_387 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_388 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_161 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_162 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_163 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_164 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_165 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_166 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_167 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_168 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_169 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_170 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_171 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_390 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_391 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_393 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_394 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_395 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_396 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_397 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_398 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_399 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_400 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_401 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_402 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_403 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_404 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_406 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_407 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_409 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_410 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_411 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_415 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_418 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_420 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_421 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_422 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_423 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_424 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_425 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_426 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_427 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_428 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_429 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_430 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_431 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_432 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_433 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_434 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_435 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_436 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_437 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_438 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_439 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_440 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_441 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_442 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_443 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_444 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_445 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_446 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_447 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_448 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_449 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_450 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_451 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_452 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_453 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_454 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_455 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_456 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_457 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_458 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_459 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_460 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_461 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_462 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_463 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_464 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_465 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_466 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_467 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_468 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_469 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_470 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_471 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_472 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_473 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_474 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_475 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_476 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_477 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_478 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_479 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_480 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_481 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_482 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_483 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_484 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_485 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_486 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_487 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_488 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_489 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_490 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_491 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_492 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_493 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_494 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_495 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_496 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_497 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_498 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_499 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_500 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_501 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_502 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_503 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_504 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_505 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_506 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_507 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_508 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_173 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_174 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_175 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_177 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_178 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_180 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_181 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_182 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_183 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_184 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_509 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_510 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_511 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_512 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_513 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_514 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_515 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_516 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_517 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_518 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_519 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_520 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_521 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_522 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_523 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_524 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_525 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_526 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_527 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_528 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_529 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_530 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_531 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_532 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_533 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_534 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_535 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_536 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_537 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_538 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_539 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_540 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_541 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_542 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_543 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_544 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_545 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_546 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_547 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_548 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_549 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_550 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_551 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_552 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_553 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_554 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_555 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_556 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_557 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_558 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_559 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_560 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_561 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_562 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_563 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_564 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_565 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_566 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_567 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_568 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_569 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_570 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_571 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_572 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_573 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_574 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_575 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_576 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_577 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_578 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_579 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_580 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_581 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_582 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_583 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_584 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_585 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_586 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_587 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_588 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_589 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_590 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_591 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_592 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_593 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_594 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_595 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_596 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_597 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_598 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_599 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_600 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_601 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_602 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_603 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_604 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_605 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_606 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_607 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_608 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_609 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_610 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_611 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_612 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_613 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_614 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_615 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_616 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_617 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_618 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_619 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_620 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_621 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_622 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_623 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_624 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_625 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_626 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_627 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_628 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_185 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_186 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_187 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_188 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_189 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_190 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_191 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_192 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_193 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_194 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_195 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_196 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_629 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_630 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_631 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_632 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_633 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_634 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_635 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_636 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_637 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_638 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_639 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_640 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_641 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_642 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_643 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_644 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_645 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_646 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_647 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_648 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_649 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_650 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_651 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_652 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_653 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_654 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_655 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_656 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_657 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_658 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_659 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_660 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_661 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_662 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_663 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_664 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_665 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_666 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_667 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_668 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_669 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_670 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_671 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_672 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_673 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_674 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_675 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_676 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_677 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_678 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_679 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_680 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_681 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_682 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_683 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_684 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_685 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_686 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_687 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_688 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_689 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_690 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_691 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_692 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_693 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_694 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_695 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_696 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_697 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_698 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_699 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_700 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_701 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_702 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_703 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_704 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_705 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_706 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_707 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_708 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_709 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_710 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_711 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_712 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_713 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_714 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_715 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_716 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_717 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_718 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_719 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_720 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_721 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_722 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_723 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_724 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_725 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_726 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_727 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_728 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_729 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_730 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_731 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_732 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_733 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_734 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_735 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_736 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_737 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_738 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_739 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_740 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_741 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_742 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_743 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_744 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_745 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_746 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_747 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_748 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_197 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_198 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_199 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_200 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_201 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_202 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_203 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_204 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_205 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_206 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_207 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_749 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_750 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_751 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_752 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_753 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_754 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_755 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_756 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_757 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_758 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_759 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_760 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_761 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_762 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_763 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_764 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_765 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_766 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_767 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_768 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_769 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_770 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_771 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_772 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_773 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_774 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_775 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_776 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_777 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_778 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_779 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_780 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_781 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_782 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_783 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_784 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_785 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_786 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_787 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_788 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_789 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_790 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_791 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_792 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_793 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_794 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_795 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_796 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_797 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_798 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_799 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_800 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_801 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_802 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_803 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_804 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_805 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_806 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_807 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_808 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_809 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_810 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_811 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_812 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_813 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_814 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_815 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_816 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_817 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_818 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_819 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_820 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_821 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_822 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_823 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_824 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_825 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_826 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_827 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_828 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_829 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_830 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_831 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_832 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_833 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_834 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_835 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_836 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_837 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_838 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_839 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_840 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_841 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_842 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_843 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_844 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_845 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_846 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_847 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_848 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_849 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_850 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_851 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_852 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_853 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_854 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_855 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_856 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_857 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_858 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_859 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_860 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_861 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_862 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_863 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_864 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_865 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_866 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_867 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_868 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_209 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_210 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_211 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_213 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_214 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_216 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_217 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_218 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_219 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_220 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_869 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_870 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_871 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_872 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_873 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_874 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_875 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_876 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_877 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_878 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_879 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_880 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_881 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_882 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_883 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_884 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_885 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_886 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_887 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_888 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_889 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_890 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_891 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_892 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_893 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_894 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_895 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_896 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_897 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_898 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_899 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_900 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_901 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_902 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_903 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_904 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_905 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_906 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_907 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_908 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_909 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_910 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_911 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_912 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_913 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_914 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_915 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_916 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_917 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_918 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_919 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_920 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_921 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_922 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_923 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_924 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_925 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_926 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_927 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_928 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_929 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_930 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_931 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_932 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_933 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_934 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_935 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_936 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_937 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_938 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_939 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_940 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_941 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_942 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_943 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_944 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_945 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_946 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_947 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_948 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_949 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_950 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_951 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_952 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_953 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_954 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_955 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_956 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_957 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_958 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_959 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_960 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_961 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_962 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_963 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_964 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_965 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_966 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_967 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_968 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_969 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_970 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_971 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_972 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_973 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_974 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_975 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_976 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_977 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_221 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_222 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_223 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_224 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_225 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_226 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_227 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_228 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_229 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_230 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_231 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_232 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_233 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_234 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_235 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_236 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_237 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_238 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_239 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_240 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_241 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_242 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_244 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_245 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_246 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_248 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_249 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_251 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_252 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_253 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_254 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_255 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_256 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_257 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_258 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_259 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_260 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_261 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_262 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_263 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_264 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_265 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_266 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_267 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_268 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1597_ (.I(\m_arbiter.o_sel_sig ),
    .Z(_1522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1598_ (.I(_1522_),
    .Z(_1523_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _1599_ (.I(_1523_),
    .ZN(_1524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1600_ (.I(_1524_),
    .Z(_1525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1601_ (.I(_1523_),
    .Z(_1526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1602_ (.I(_1526_),
    .Z(_1527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1603_ (.A1(_1527_),
    .A2(\m_arbiter.wb0_o_dat[7] ),
    .Z(_1528_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1604_ (.A1(_1525_),
    .A2(net41),
    .B(_1528_),
    .ZN(_1529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1605_ (.I(net237),
    .ZN(net147),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1606_ (.A1(_1527_),
    .A2(\m_arbiter.wb0_o_dat[6] ),
    .Z(_1530_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1607_ (.A1(_1525_),
    .A2(net40),
    .B(_1530_),
    .ZN(_1531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1608_ (.I(net236),
    .ZN(net146),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1609_ (.A1(_1527_),
    .A2(\m_arbiter.wb0_o_dat[5] ),
    .Z(_1532_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1610_ (.A1(_1525_),
    .A2(net39),
    .B(_1532_),
    .ZN(_1533_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1611_ (.I(net235),
    .ZN(net145),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1612_ (.A1(_1527_),
    .A2(\m_arbiter.wb0_o_dat[4] ),
    .Z(_1534_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1613_ (.A1(_1525_),
    .A2(net38),
    .B(_1534_),
    .ZN(_1535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1614_ (.I(net234),
    .ZN(net144),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1615_ (.A1(_1527_),
    .A2(net37),
    .ZN(_1536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1616_ (.A1(_1525_),
    .A2(\m_arbiter.wb0_o_dat[3] ),
    .ZN(_1537_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1617_ (.A1(_1536_),
    .A2(_1537_),
    .Z(_1538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1618_ (.I(_1538_),
    .Z(_1539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1619_ (.I(_1539_),
    .ZN(net143),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _1620_ (.I(_1526_),
    .Z(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1621_ (.A1(_1540_),
    .A2(net36),
    .ZN(_1541_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1622_ (.A1(_1524_),
    .A2(\m_arbiter.wb0_o_dat[2] ),
    .ZN(_1542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1623_ (.A1(_1541_),
    .A2(_1542_),
    .Z(_1543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1624_ (.I(_1543_),
    .Z(_1544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1625_ (.I(_1544_),
    .ZN(net142),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1626_ (.A1(_1540_),
    .A2(net35),
    .ZN(_1545_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1627_ (.A1(_1524_),
    .A2(\m_arbiter.wb0_o_dat[1] ),
    .ZN(_1546_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1628_ (.A1(_1545_),
    .A2(_1546_),
    .Z(_1547_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1629_ (.I(_1547_),
    .Z(_1548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1630_ (.I(_1548_),
    .ZN(net141),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1631_ (.A1(_1527_),
    .A2(net28),
    .ZN(_1549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1632_ (.A1(_1525_),
    .A2(net531),
    .ZN(_1550_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1633_ (.A1(_1549_),
    .A2(_1550_),
    .Z(_1551_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1634_ (.I(_1551_),
    .Z(_1552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1635_ (.I(_1552_),
    .ZN(net134),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1636_ (.I(net490),
    .Z(_1553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1637_ (.I(_1553_),
    .Z(_1554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1638_ (.I(\m_arbiter.wb0_adr[8] ),
    .ZN(_1555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1639_ (.A1(_1523_),
    .A2(net25),
    .ZN(_1556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _1640_ (.I(_1522_),
    .Z(_1557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _1641_ (.I0(\m_arbiter.wb0_adr[9] ),
    .I1(net26),
    .S(_1557_),
    .Z(_1558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1642_ (.A1(_1526_),
    .A2(_1555_),
    .B(_1556_),
    .C(_1558_),
    .ZN(_1559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1643_ (.I0(\m_arbiter.wb0_adr[14] ),
    .I1(net8),
    .S(net389),
    .Z(_1560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1644_ (.I0(\m_arbiter.wb0_adr[15] ),
    .I1(net9),
    .S(_1522_),
    .Z(_1561_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1645_ (.A1(_1560_),
    .A2(_1561_),
    .ZN(_1562_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1646_ (.I0(\m_arbiter.wb0_adr[7] ),
    .I1(net24),
    .S(_1557_),
    .Z(_1563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1647_ (.I0(\m_arbiter.wb0_adr[6] ),
    .I1(net23),
    .S(_1523_),
    .Z(_1564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1648_ (.A1(_1563_),
    .A2(_1564_),
    .Z(_1565_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1649_ (.I(net90),
    .ZN(_1566_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1650_ (.I0(\m_arbiter.wb0_adr[13] ),
    .I1(net7),
    .S(_1522_),
    .Z(_1567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1651_ (.A1(_1566_),
    .A2(_1567_),
    .ZN(_1568_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1652_ (.A1(_1559_),
    .A2(_1562_),
    .A3(_1565_),
    .A4(_1568_),
    .ZN(_1569_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _1653_ (.I0(\m_arbiter.wb0_adr[12] ),
    .I1(net6),
    .S(_1523_),
    .Z(_1570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1654_ (.I0(\m_arbiter.wb0_adr[22] ),
    .I1(net17),
    .S(_1523_),
    .Z(_1571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1655_ (.I0(\m_arbiter.wb0_adr[21] ),
    .I1(net16),
    .S(_1523_),
    .Z(_1572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1656_ (.A1(_1570_),
    .A2(_1571_),
    .A3(_1572_),
    .ZN(_1573_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1657_ (.I0(\m_arbiter.wb0_adr[16] ),
    .I1(net10),
    .S(_1557_),
    .Z(_1574_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1658_ (.I0(\m_arbiter.wb0_adr[18] ),
    .I1(net12),
    .S(_1557_),
    .Z(_1575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1659_ (.A1(_1574_),
    .A2(_1575_),
    .ZN(_1576_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1660_ (.I(\m_arbiter.wb0_adr[23] ),
    .ZN(_1577_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1661_ (.A1(_1526_),
    .A2(net18),
    .ZN(_1578_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _1662_ (.I0(\m_arbiter.wb0_adr[20] ),
    .I1(net15),
    .S(_1523_),
    .Z(_1579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1663_ (.A1(_1526_),
    .A2(_1577_),
    .B(_1578_),
    .C(_1579_),
    .ZN(_1580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _1664_ (.I0(\m_arbiter.wb0_adr[11] ),
    .I1(net5),
    .S(_1557_),
    .Z(_1581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1665_ (.I0(\m_arbiter.wb0_adr[10] ),
    .I1(net4),
    .S(_1557_),
    .Z(_1582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1666_ (.I0(\m_arbiter.wb0_adr[19] ),
    .I1(net13),
    .S(_1557_),
    .Z(_1583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1667_ (.I0(\m_arbiter.wb0_adr[17] ),
    .I1(net11),
    .S(_1557_),
    .Z(_1584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1668_ (.A1(_1581_),
    .A2(_1582_),
    .A3(_1583_),
    .A4(_1584_),
    .ZN(_1585_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1669_ (.A1(_1573_),
    .A2(_1576_),
    .A3(_1580_),
    .A4(_1585_),
    .ZN(_1586_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1670_ (.A1(_1569_),
    .A2(_1586_),
    .B(net90),
    .ZN(_1587_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1671_ (.I0(\m_arbiter.wb0_adr[1] ),
    .I1(net14),
    .S(net388),
    .Z(_1588_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1672_ (.I(_1588_),
    .Z(net128),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1673_ (.I0(\m_arbiter.wb0_adr[0] ),
    .I1(net3),
    .S(_1523_),
    .Z(_1589_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1674_ (.I(_1589_),
    .Z(net127),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1675_ (.A1(net128),
    .A2(net127),
    .ZN(_1590_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1676_ (.I0(\m_arbiter.wb0_adr[5] ),
    .I1(net22),
    .S(_1557_),
    .Z(_1591_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1677_ (.I(_1591_),
    .Z(net132),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1678_ (.I0(\m_arbiter.wb0_adr[4] ),
    .I1(net21),
    .S(_1522_),
    .Z(_1592_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1679_ (.I(_1592_),
    .Z(net131),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _1680_ (.I(net131),
    .ZN(_1593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1681_ (.A1(_1565_),
    .A2(net132),
    .A3(_1593_),
    .ZN(_1594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1682_ (.A1(_1574_),
    .A2(_1575_),
    .A3(_1583_),
    .A4(_1584_),
    .ZN(_0390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1683_ (.I0(\m_arbiter.wb0_adr[23] ),
    .I1(net18),
    .S(_1523_),
    .Z(_0391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1684_ (.A1(_0391_),
    .A2(_1579_),
    .ZN(_0392_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1685_ (.A1(_1571_),
    .A2(_1572_),
    .ZN(_0393_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1686_ (.A1(_0390_),
    .A2(_0392_),
    .A3(_0393_),
    .Z(_0394_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1687_ (.A1(_1560_),
    .A2(_1561_),
    .A3(_1567_),
    .ZN(_0395_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1688_ (.I0(\m_arbiter.wb0_adr[8] ),
    .I1(net25),
    .S(_1557_),
    .Z(_0396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1689_ (.A1(_0396_),
    .A2(_1558_),
    .A3(_1581_),
    .A4(_1582_),
    .ZN(_0397_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1690_ (.I0(\m_arbiter.wb0_adr[3] ),
    .I1(net20),
    .S(_1522_),
    .Z(_0398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1691_ (.I(_0398_),
    .Z(net130),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1692_ (.I0(\m_arbiter.wb0_adr[2] ),
    .I1(net19),
    .S(net388),
    .Z(_0399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1693_ (.I(_0399_),
    .Z(net129),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1694_ (.A1(net130),
    .A2(net129),
    .ZN(_0400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1695_ (.A1(_1570_),
    .A2(net255),
    .A3(net247),
    .A4(_0400_),
    .Z(_0401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1696_ (.A1(_1590_),
    .A2(_1594_),
    .A3(_0394_),
    .A4(_0401_),
    .ZN(_0402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1697_ (.A1(net248),
    .A2(_0392_),
    .A3(_0393_),
    .ZN(_0403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1698_ (.A1(_1570_),
    .A2(net255),
    .A3(net246),
    .A4(_0400_),
    .ZN(_0404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1699_ (.A1(_1563_),
    .A2(_1564_),
    .ZN(_0405_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _1700_ (.I(net132),
    .ZN(_0406_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1701_ (.A1(_0405_),
    .A2(_0406_),
    .A3(_1593_),
    .ZN(_0407_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1702_ (.I(net128),
    .ZN(_0408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1703_ (.A1(_0408_),
    .A2(net127),
    .ZN(_0409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _1704_ (.A1(_0403_),
    .A2(_0404_),
    .A3(_0407_),
    .A4(_0409_),
    .Z(_0410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1705_ (.A1(_1587_),
    .A2(_0402_),
    .A3(_0410_),
    .Z(_0411_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _1706_ (.I(_0411_),
    .Z(_0412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1707_ (.I(_0412_),
    .Z(_0413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1708_ (.I(\wb_cross_clk.m_wb_i_dat[15] ),
    .ZN(_0414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1709_ (.I(_1553_),
    .Z(_0415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1710_ (.A1(_0414_),
    .A2(_0415_),
    .ZN(_0416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1711_ (.A1(_1554_),
    .A2(\wb_compressor.wb_i_dat[15] ),
    .B(_0413_),
    .C(_0416_),
    .ZN(_0417_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1712_ (.A1(net255),
    .A2(net247),
    .ZN(_0418_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1713_ (.A1(_0391_),
    .A2(_1579_),
    .ZN(_0419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1714_ (.A1(_0405_),
    .A2(_0393_),
    .A3(_0419_),
    .ZN(_0420_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1715_ (.A1(_1566_),
    .A2(_1570_),
    .ZN(_0421_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1716_ (.A1(_0391_),
    .A2(_1579_),
    .B(_0390_),
    .C(_0421_),
    .ZN(_0422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1717_ (.A1(_1573_),
    .A2(_1576_),
    .A3(_1580_),
    .A4(_1585_),
    .Z(_0423_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1718_ (.A1(_1559_),
    .A2(_1562_),
    .A3(_1565_),
    .A4(_1568_),
    .Z(_0424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1719_ (.A1(_0418_),
    .A2(_0420_),
    .A3(_0422_),
    .B1(_0423_),
    .B2(_0424_),
    .ZN(_0425_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1720_ (.I(_0425_),
    .Z(_0426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1721_ (.A1(\iram_latched[15] ),
    .A2(_0426_),
    .ZN(_0427_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1722_ (.A1(_0417_),
    .A2(_0427_),
    .ZN(net117),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1723_ (.I(_1553_),
    .Z(_0428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1724_ (.I(\wb_cross_clk.m_wb_i_dat[14] ),
    .ZN(_0429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1725_ (.A1(_0429_),
    .A2(_0415_),
    .ZN(_0430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1726_ (.A1(_0428_),
    .A2(\wb_compressor.wb_i_dat[14] ),
    .B(_0413_),
    .C(_0430_),
    .ZN(_0431_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1727_ (.A1(\iram_latched[14] ),
    .A2(_0426_),
    .ZN(_0432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1728_ (.A1(_0431_),
    .A2(_0432_),
    .ZN(net116),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1729_ (.I(\wb_cross_clk.m_wb_i_dat[13] ),
    .ZN(_0433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1730_ (.A1(_0433_),
    .A2(_0415_),
    .ZN(_0434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1731_ (.A1(_0428_),
    .A2(\wb_compressor.wb_i_dat[13] ),
    .B(_0412_),
    .C(_0434_),
    .ZN(_0435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1732_ (.A1(\iram_latched[13] ),
    .A2(_0426_),
    .ZN(_0436_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1733_ (.A1(_0435_),
    .A2(_0436_),
    .ZN(net115),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1734_ (.I(\wb_cross_clk.m_wb_i_dat[12] ),
    .ZN(_0437_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1735_ (.A1(_0437_),
    .A2(_0415_),
    .ZN(_0438_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1736_ (.A1(_0428_),
    .A2(\wb_compressor.wb_i_dat[12] ),
    .B(_0412_),
    .C(_0438_),
    .ZN(_0439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1737_ (.A1(\iram_latched[12] ),
    .A2(_0426_),
    .ZN(_0440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1738_ (.A1(_0439_),
    .A2(_0440_),
    .ZN(net114),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1739_ (.I(\wb_cross_clk.m_wb_i_dat[11] ),
    .ZN(_0441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1740_ (.A1(_0441_),
    .A2(_0415_),
    .ZN(_0442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1741_ (.A1(_0428_),
    .A2(\wb_compressor.wb_i_dat[11] ),
    .B(_0412_),
    .C(_0442_),
    .ZN(_0443_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1742_ (.A1(\iram_latched[11] ),
    .A2(_0426_),
    .ZN(_0444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1743_ (.A1(_0443_),
    .A2(_0444_),
    .ZN(net113),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1744_ (.I(\wb_cross_clk.m_wb_i_dat[10] ),
    .ZN(_0445_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1745_ (.A1(_0445_),
    .A2(_0415_),
    .ZN(_0446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1746_ (.A1(_0428_),
    .A2(\wb_compressor.wb_i_dat[10] ),
    .B(_0412_),
    .C(_0446_),
    .ZN(_0447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1747_ (.A1(\iram_latched[10] ),
    .A2(_0426_),
    .ZN(_0448_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1748_ (.A1(_0447_),
    .A2(_0448_),
    .ZN(net112),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1749_ (.I(\wb_cross_clk.m_wb_i_dat[9] ),
    .ZN(_0449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1750_ (.A1(_0449_),
    .A2(_0415_),
    .ZN(_0450_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1751_ (.A1(_0428_),
    .A2(\wb_compressor.wb_i_dat[9] ),
    .B(_0412_),
    .C(_0450_),
    .ZN(_0451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1752_ (.A1(\iram_latched[9] ),
    .A2(_0426_),
    .ZN(_0452_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1753_ (.A1(_0451_),
    .A2(_0452_),
    .ZN(net126),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1754_ (.I(\wb_cross_clk.m_wb_i_dat[8] ),
    .ZN(_0453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1755_ (.A1(_0453_),
    .A2(_0415_),
    .ZN(_0454_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1756_ (.A1(_0428_),
    .A2(\wb_compressor.wb_i_dat[8] ),
    .B(_0412_),
    .C(_0454_),
    .ZN(_0455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1757_ (.A1(\iram_latched[8] ),
    .A2(_0426_),
    .ZN(_0456_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1758_ (.A1(_0455_),
    .A2(_0456_),
    .ZN(net125),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1759_ (.I(_0426_),
    .Z(_0457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _1760_ (.I(_1553_),
    .Z(_0458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1761_ (.I0(\wb_compressor.wb_i_dat[7] ),
    .I1(\wb_cross_clk.m_wb_i_dat[7] ),
    .S(_0458_),
    .Z(_0459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1762_ (.A1(\iram_latched[7] ),
    .A2(_0457_),
    .B1(_0459_),
    .B2(_0413_),
    .ZN(_0460_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1763_ (.A1(_1590_),
    .A2(_1594_),
    .A3(_0394_),
    .A4(_0401_),
    .Z(_0461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1764_ (.I(_0461_),
    .Z(_0462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1765_ (.I(net127),
    .ZN(_0463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1766_ (.A1(net128),
    .A2(_0463_),
    .ZN(_0464_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1767_ (.A1(net128),
    .A2(_0463_),
    .ZN(_0465_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1768_ (.I(_0465_),
    .ZN(_0466_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1769_ (.A1(_1526_),
    .A2(\m_arbiter.wb0_adr[12] ),
    .Z(_0467_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1770_ (.A1(_1524_),
    .A2(net6),
    .B(_0467_),
    .ZN(_0468_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1771_ (.A1(net130),
    .A2(net129),
    .Z(_0469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1772_ (.A1(_0468_),
    .A2(_0403_),
    .A3(_0418_),
    .A4(_0469_),
    .ZN(_0470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1773_ (.A1(_0464_),
    .A2(_0466_),
    .B(net231),
    .C(net241),
    .ZN(_0471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1774_ (.A1(net97),
    .A2(_0471_),
    .ZN(_0472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1775_ (.A1(_0405_),
    .A2(_0406_),
    .A3(net131),
    .ZN(_0473_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1776_ (.A1(_0473_),
    .A2(_0403_),
    .A3(_0404_),
    .A4(_0465_),
    .ZN(_0474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1777_ (.A1(_0473_),
    .A2(_0403_),
    .A3(_0404_),
    .A4(_0409_),
    .ZN(_0475_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1778_ (.A1(net174),
    .A2(net228),
    .B1(net224),
    .B2(net201),
    .ZN(_0476_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1779_ (.A1(_0472_),
    .A2(_0476_),
    .ZN(_0477_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1780_ (.A1(_0462_),
    .A2(_0477_),
    .ZN(_0478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1781_ (.A1(_0460_),
    .A2(_0478_),
    .ZN(net124),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1782_ (.I0(\wb_compressor.wb_i_dat[6] ),
    .I1(\wb_cross_clk.m_wb_i_dat[6] ),
    .S(_0458_),
    .Z(_0479_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1783_ (.A1(\iram_latched[6] ),
    .A2(_0457_),
    .B1(_0479_),
    .B2(_0413_),
    .ZN(_0480_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1784_ (.A1(net96),
    .A2(_0471_),
    .ZN(_0481_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1785_ (.A1(net173),
    .A2(net227),
    .B1(net223),
    .B2(net200),
    .ZN(_0482_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1786_ (.A1(_0481_),
    .A2(_0482_),
    .ZN(_0483_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1787_ (.A1(_0462_),
    .A2(_0483_),
    .ZN(_0484_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1788_ (.A1(_0480_),
    .A2(_0484_),
    .ZN(net123),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1789_ (.I0(\wb_compressor.wb_i_dat[5] ),
    .I1(\wb_cross_clk.m_wb_i_dat[5] ),
    .S(_0458_),
    .Z(_0485_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1790_ (.A1(\iram_latched[5] ),
    .A2(_0457_),
    .B1(_0485_),
    .B2(_0413_),
    .ZN(_0486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1791_ (.A1(net95),
    .A2(_0471_),
    .ZN(_0487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1792_ (.A1(net172),
    .A2(net227),
    .B1(net223),
    .B2(net199),
    .ZN(_0488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1793_ (.A1(_0487_),
    .A2(_0488_),
    .ZN(_0489_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1794_ (.A1(_0462_),
    .A2(_0489_),
    .ZN(_0490_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1795_ (.A1(_0486_),
    .A2(_0490_),
    .ZN(net122),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1796_ (.I0(\wb_compressor.wb_i_dat[4] ),
    .I1(\wb_cross_clk.m_wb_i_dat[4] ),
    .S(_0458_),
    .Z(_0491_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1797_ (.A1(\iram_latched[4] ),
    .A2(_0457_),
    .B1(_0491_),
    .B2(_0413_),
    .ZN(_0492_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1798_ (.A1(net94),
    .A2(_0471_),
    .ZN(_0493_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1799_ (.A1(net171),
    .A2(net226),
    .B1(net222),
    .B2(net198),
    .ZN(_0494_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1800_ (.A1(_0493_),
    .A2(_0494_),
    .ZN(_0495_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1801_ (.A1(_0462_),
    .A2(_0495_),
    .ZN(_0496_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1802_ (.A1(_0492_),
    .A2(_0496_),
    .ZN(net121),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1803_ (.I0(\wb_compressor.wb_i_dat[3] ),
    .I1(\wb_cross_clk.m_wb_i_dat[3] ),
    .S(_0458_),
    .Z(_0497_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1804_ (.A1(\iram_latched[3] ),
    .A2(_0457_),
    .B1(_0497_),
    .B2(_0413_),
    .ZN(_0498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1805_ (.A1(net93),
    .A2(_0471_),
    .ZN(_0499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1806_ (.A1(net170),
    .A2(net226),
    .B1(net222),
    .B2(net197),
    .ZN(_0500_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1807_ (.A1(_0499_),
    .A2(_0500_),
    .ZN(_0501_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1808_ (.A1(_0462_),
    .A2(_0501_),
    .ZN(_0502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1809_ (.A1(_0498_),
    .A2(_0502_),
    .ZN(net120),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1810_ (.I0(\wb_compressor.wb_i_dat[2] ),
    .I1(\wb_cross_clk.m_wb_i_dat[2] ),
    .S(_0458_),
    .Z(_0503_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1811_ (.A1(\iram_latched[2] ),
    .A2(_0457_),
    .B1(_0503_),
    .B2(_0413_),
    .ZN(_0504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1812_ (.A1(net86),
    .A2(_0471_),
    .ZN(_0505_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1813_ (.A1(net169),
    .A2(net225),
    .B1(net221),
    .B2(net194),
    .ZN(_0506_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1814_ (.A1(_0505_),
    .A2(_0506_),
    .ZN(_0507_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1815_ (.A1(_0462_),
    .A2(_0507_),
    .ZN(_0508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1816_ (.A1(_0504_),
    .A2(_0508_),
    .ZN(net119),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1817_ (.I0(\wb_compressor.wb_i_dat[1] ),
    .I1(\wb_cross_clk.m_wb_i_dat[1] ),
    .S(_0458_),
    .Z(_0509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1818_ (.A1(\iram_latched[1] ),
    .A2(_0457_),
    .B1(_0509_),
    .B2(_0413_),
    .ZN(_0510_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1819_ (.A1(net77),
    .A2(_0471_),
    .ZN(_0511_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1820_ (.A1(net162),
    .A2(net225),
    .B1(net221),
    .B2(net186),
    .ZN(_0512_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1821_ (.A1(_0512_),
    .A2(_0511_),
    .ZN(_0513_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1822_ (.A1(_0462_),
    .A2(_0513_),
    .ZN(_0514_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1823_ (.A1(_0510_),
    .A2(_0514_),
    .ZN(net118),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1824_ (.I0(\wb_compressor.wb_i_dat[0] ),
    .I1(\wb_cross_clk.m_wb_i_dat[0] ),
    .S(_0415_),
    .Z(_0515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1825_ (.A1(\iram_latched[0] ),
    .A2(_0457_),
    .B1(_0515_),
    .B2(_0413_),
    .ZN(_0516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1826_ (.A1(net66),
    .A2(_0471_),
    .ZN(_0517_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1827_ (.A1(net151),
    .A2(net225),
    .B1(net221),
    .B2(net175),
    .ZN(_0518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1828_ (.A1(_0518_),
    .A2(_0517_),
    .ZN(_0519_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1829_ (.A1(_0462_),
    .A2(_0519_),
    .ZN(_0520_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1830_ (.A1(_0520_),
    .A2(_0516_),
    .ZN(net111),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1831_ (.I(\wb_compressor.wb_ack ),
    .ZN(_0521_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1832_ (.A1(_1524_),
    .A2(\m_arbiter.i_wb0_cyc ),
    .ZN(_0522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1833_ (.A1(_1526_),
    .A2(net27),
    .ZN(_0523_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1834_ (.I(net108),
    .Z(_0524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1835_ (.A1(_0522_),
    .A2(_0523_),
    .B(_0524_),
    .ZN(_0525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1836_ (.A1(_1524_),
    .A2(net46),
    .Z(_0526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1837_ (.A1(_0525_),
    .A2(_0526_),
    .ZN(_0527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1838_ (.I(\wb_cross_clk.ack_next_hold ),
    .ZN(_0528_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1839_ (.A1(_0528_),
    .A2(\wb_cross_clk.m_s_sync.d_data[46] ),
    .A3(net490),
    .ZN(_0529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1840_ (.A1(_1553_),
    .A2(_0527_),
    .B(_0529_),
    .ZN(_0530_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1841_ (.A1(_0521_),
    .A2(_0412_),
    .A3(net491),
    .ZN(_0531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1842_ (.A1(\wb_compressor.state[6] ),
    .A2(_0531_),
    .ZN(_0532_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1843_ (.A1(net85),
    .A2(net84),
    .B(_0411_),
    .C(_0530_),
    .ZN(_0533_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1844_ (.I(_0533_),
    .ZN(_0534_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1845_ (.I(\wb_compressor.burst_end[0] ),
    .ZN(_0535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1846_ (.A1(\wb_compressor.burst_cnt[0] ),
    .A2(\wb_compressor.burst_cnt[1] ),
    .Z(_0536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1847_ (.A1(\wb_compressor.burst_cnt[0] ),
    .A2(\wb_compressor.burst_cnt[1] ),
    .ZN(_0537_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1848_ (.A1(\wb_compressor.burst_end[0] ),
    .A2(_0537_),
    .Z(_0538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1849_ (.A1(\wb_compressor.burst_end[2] ),
    .A2(\wb_compressor.burst_cnt[2] ),
    .ZN(_0539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1850_ (.A1(_0535_),
    .A2(_0536_),
    .B(_0538_),
    .C(_0539_),
    .ZN(_0540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1851_ (.A1(\wb_compressor.state[4] ),
    .A2(_0534_),
    .A3(_0540_),
    .ZN(_0541_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1852_ (.I(net193),
    .Z(_0542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1853_ (.I(_0542_),
    .Z(_0543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1854_ (.I(_0543_),
    .Z(_0544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1855_ (.A1(_0532_),
    .A2(_0541_),
    .B(_0544_),
    .ZN(_0014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1856_ (.A1(_0533_),
    .A2(_0540_),
    .B(\wb_compressor.state[5] ),
    .ZN(_0545_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1857_ (.I(\wb_compressor.l_we ),
    .ZN(_0546_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1858_ (.A1(net84),
    .A2(\wb_compressor.state[2] ),
    .Z(_0547_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1859_ (.A1(_0546_),
    .A2(_0547_),
    .ZN(_0548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1860_ (.A1(_0545_),
    .A2(_0548_),
    .B(_0544_),
    .ZN(_0013_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1861_ (.I(_0543_),
    .Z(_0549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1862_ (.I(\wb_compressor.state[6] ),
    .ZN(_0550_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1863_ (.A1(_0550_),
    .A2(_0531_),
    .ZN(_0551_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1864_ (.A1(\wb_compressor.state[4] ),
    .A2(_0533_),
    .B1(_0547_),
    .B2(\wb_compressor.l_we ),
    .C(_0551_),
    .ZN(_0552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1865_ (.A1(_0549_),
    .A2(net205),
    .ZN(_0012_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1866_ (.I(_0542_),
    .Z(_0553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1867_ (.I(net84),
    .ZN(_0554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1868_ (.I(\wb_compressor.state[3] ),
    .Z(_0555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1869_ (.I(_0555_),
    .Z(_0556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1870_ (.A1(_0554_),
    .A2(\wb_compressor.state[2] ),
    .B(_0556_),
    .ZN(_0557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1871_ (.A1(_0553_),
    .A2(_0557_),
    .ZN(_0011_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _1872_ (.I(net490),
    .ZN(_0558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _1873_ (.I(_0558_),
    .Z(_0559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1874_ (.I0(\wb_cross_clk.m_s_sync.d_data[41] ),
    .I1(_1583_),
    .S(_0559_),
    .Z(_0560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1875_ (.I0(\wb_cross_clk.m_s_sync.d_data[35] ),
    .I1(net507),
    .S(_0559_),
    .Z(_0561_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1876_ (.I0(\wb_cross_clk.m_s_sync.d_data[37] ),
    .I1(net524),
    .S(_0559_),
    .Z(_0562_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1877_ (.A1(_0560_),
    .A2(_0561_),
    .A3(_0562_),
    .ZN(_0563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1878_ (.I0(\wb_cross_clk.m_s_sync.d_data[38] ),
    .I1(_1574_),
    .S(_0559_),
    .Z(_0564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1879_ (.I0(\wb_cross_clk.m_s_sync.d_data[42] ),
    .I1(_1579_),
    .S(_0558_),
    .Z(_0565_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1880_ (.I0(\wb_cross_clk.m_s_sync.d_data[40] ),
    .I1(_1575_),
    .S(_0558_),
    .Z(_0566_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1881_ (.I0(\wb_cross_clk.m_s_sync.d_data[45] ),
    .I1(_0391_),
    .S(_0559_),
    .Z(_0567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1882_ (.A1(_0564_),
    .A2(_0565_),
    .A3(_0566_),
    .A4(_0567_),
    .ZN(_0568_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1883_ (.I0(\wb_cross_clk.m_s_sync.d_data[39] ),
    .I1(_1584_),
    .S(_0558_),
    .Z(_0569_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1884_ (.I0(\wb_cross_clk.m_s_sync.d_data[36] ),
    .I1(net518),
    .S(_0558_),
    .Z(_0570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1885_ (.I0(\wb_cross_clk.m_s_sync.d_data[44] ),
    .I1(_1571_),
    .S(_0558_),
    .Z(_0571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1886_ (.I0(\wb_cross_clk.m_s_sync.d_data[43] ),
    .I1(net521),
    .S(_0559_),
    .Z(_0572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1887_ (.A1(_0569_),
    .A2(_0570_),
    .A3(_0571_),
    .A4(_0572_),
    .ZN(_0573_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1888_ (.A1(_0563_),
    .A2(_0568_),
    .A3(_0573_),
    .ZN(_0574_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1889_ (.A1(_0411_),
    .A2(net491),
    .A3(_0574_),
    .ZN(_0575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1890_ (.A1(\wb_compressor.state[0] ),
    .A2(_0575_),
    .ZN(_0576_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1891_ (.A1(\wb_compressor.state[1] ),
    .A2(_0542_),
    .ZN(_0577_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1892_ (.A1(_0576_),
    .A2(_0577_),
    .ZN(_0010_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1893_ (.I(\sspi.state[1] ),
    .ZN(_0578_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1894_ (.I(_0524_),
    .Z(_0579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1895_ (.I(_0579_),
    .Z(_0580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1896_ (.I(\sspi.sy_clk[2] ),
    .ZN(_0581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1897_ (.A1(_0581_),
    .A2(\sspi.sy_clk[3] ),
    .ZN(_0582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1898_ (.A1(_0426_),
    .A2(_0527_),
    .ZN(_0583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1899_ (.A1(\wb_cross_clk.msy_xor_err ),
    .A2(\wb_cross_clk.prev_xor_err ),
    .ZN(_0584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1900_ (.A1(_1553_),
    .A2(net262),
    .ZN(_0585_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1901_ (.A1(\wb_compressor.wb_err ),
    .A2(_1553_),
    .B(_0585_),
    .ZN(_0586_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1902_ (.A1(_1587_),
    .A2(_0402_),
    .A3(_0410_),
    .A4(_0586_),
    .ZN(_0587_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1903_ (.A1(_0403_),
    .A2(net500),
    .A3(_0407_),
    .A4(_0409_),
    .ZN(_0588_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1904_ (.A1(_0462_),
    .A2(_0588_),
    .ZN(_0589_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1905_ (.A1(_1587_),
    .A2(_0583_),
    .B(_0587_),
    .C(net219),
    .ZN(_0590_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1906_ (.A1(_0525_),
    .A2(_0526_),
    .Z(_0591_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1907_ (.A1(iram_wb_ack_del),
    .A2(net229),
    .B1(_0591_),
    .B2(_0462_),
    .C(_0588_),
    .ZN(_0592_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1908_ (.A1(\wb_cross_clk.msy_xor_ack ),
    .A2(\wb_cross_clk.prev_xor_ack ),
    .ZN(_0593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1909_ (.A1(_1553_),
    .A2(net260),
    .ZN(_0594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1910_ (.A1(\wb_compressor.wb_ack ),
    .A2(_1553_),
    .B(_0594_),
    .ZN(_0595_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1911_ (.I0(net218),
    .I1(_0595_),
    .S(_0412_),
    .Z(_0596_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1912_ (.A1(_0590_),
    .A2(_0596_),
    .B(_0522_),
    .ZN(_0597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1913_ (.A1(_0582_),
    .A2(_0597_),
    .ZN(_0598_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1914_ (.A1(_0524_),
    .A2(_0582_),
    .ZN(_0599_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1915_ (.I(\sspi.bit_cnt[4] ),
    .ZN(_0600_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _1916_ (.I(\sspi.bit_cnt[1] ),
    .ZN(_0601_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _1917_ (.I(\sspi.bit_cnt[0] ),
    .ZN(_0602_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1918_ (.A1(_0601_),
    .A2(_0602_),
    .ZN(_0603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1919_ (.A1(\sspi.bit_cnt[1] ),
    .A2(\sspi.bit_cnt[0] ),
    .ZN(_0604_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1920_ (.A1(\sspi.bit_cnt[2] ),
    .A2(net259),
    .Z(_0605_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1921_ (.A1(_0603_),
    .A2(_0605_),
    .ZN(_0606_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1922_ (.A1(_0601_),
    .A2(_0602_),
    .ZN(_0607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1923_ (.A1(\sspi.bit_cnt[2] ),
    .A2(_0607_),
    .B(\sspi.bit_cnt[3] ),
    .ZN(_0608_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _1924_ (.I(\sspi.bit_cnt[3] ),
    .ZN(_0609_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _1925_ (.I(\sspi.bit_cnt[2] ),
    .ZN(_0610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1926_ (.A1(_0609_),
    .A2(_0610_),
    .A3(net259),
    .ZN(_0611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1927_ (.A1(_0608_),
    .A2(_0611_),
    .Z(_0612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1928_ (.A1(_0606_),
    .A2(_0612_),
    .ZN(_0613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1929_ (.A1(_0600_),
    .A2(_0582_),
    .A3(_0613_),
    .ZN(_0614_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1930_ (.A1(_0524_),
    .A2(_0614_),
    .ZN(_0615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1931_ (.A1(\sspi.state[5] ),
    .A2(_0599_),
    .B1(_0615_),
    .B2(\sspi.state[7] ),
    .ZN(_0616_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1932_ (.A1(_0578_),
    .A2(_0580_),
    .A3(_0598_),
    .B(_0616_),
    .ZN(_0007_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1933_ (.I(\sspi.state[5] ),
    .ZN(_0617_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1934_ (.A1(_0581_),
    .A2(\sspi.sy_clk[3] ),
    .Z(_0618_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1935_ (.I(net92),
    .Z(_0619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1936_ (.A1(_0619_),
    .A2(_0618_),
    .ZN(_0620_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1937_ (.I(\sspi.state[0] ),
    .ZN(_0621_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _1938_ (.I(_0524_),
    .ZN(_0622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1939_ (.I(_0622_),
    .Z(_0623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1940_ (.A1(_0617_),
    .A2(_0618_),
    .B1(_0620_),
    .B2(_0621_),
    .C(_0623_),
    .ZN(_0002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1941_ (.I(\sspi.state[3] ),
    .ZN(_0624_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1942_ (.A1(\sspi.state[7] ),
    .A2(_0614_),
    .ZN(_0625_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1943_ (.A1(_0624_),
    .A2(_0598_),
    .B(_0625_),
    .ZN(_0626_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1944_ (.A1(_0623_),
    .A2(_0626_),
    .Z(_0627_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1945_ (.I(_0627_),
    .Z(_0009_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1946_ (.A1(\sspi.state[6] ),
    .A2(_0614_),
    .ZN(_0628_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1947_ (.I(_0619_),
    .Z(_0629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1948_ (.A1(\sspi.state[2] ),
    .A2(_0629_),
    .A3(_0582_),
    .ZN(_0630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1949_ (.I(_0579_),
    .Z(_0631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1950_ (.A1(_0628_),
    .A2(_0630_),
    .B(_0631_),
    .ZN(_0008_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1951_ (.A1(_0622_),
    .A2(_0598_),
    .ZN(_0632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1952_ (.A1(\sspi.state[6] ),
    .A2(_0615_),
    .ZN(_0633_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1953_ (.A1(_0578_),
    .A2(_0632_),
    .B(_0633_),
    .ZN(_0003_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1954_ (.I(_0579_),
    .Z(_0634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1955_ (.A1(_0608_),
    .A2(_0611_),
    .ZN(_0635_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1956_ (.I(_0635_),
    .Z(_0636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1957_ (.A1(_0600_),
    .A2(_0606_),
    .A3(_0636_),
    .ZN(_0637_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1958_ (.A1(_0582_),
    .A2(net230),
    .ZN(_0638_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1959_ (.I(\sspi.state[4] ),
    .Z(_0639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1960_ (.A1(\sspi.state[0] ),
    .A2(_0620_),
    .B1(_0638_),
    .B2(_0639_),
    .ZN(_0640_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1961_ (.A1(_0634_),
    .A2(_0640_),
    .ZN(_0006_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1962_ (.I(_0622_),
    .Z(_0641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1963_ (.A1(_0641_),
    .A2(\sspi.state[2] ),
    .A3(_0620_),
    .ZN(_0642_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1964_ (.A1(_0624_),
    .A2(_0632_),
    .B(_0642_),
    .ZN(_0005_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1965_ (.A1(_0641_),
    .A2(_0639_),
    .ZN(_0643_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1966_ (.A1(\sspi.state[2] ),
    .A2(_0599_),
    .ZN(_0644_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1967_ (.A1(_0638_),
    .A2(_0643_),
    .B(_0644_),
    .ZN(_0004_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1968_ (.I0(\m_arbiter.wb0_o_dat[8] ),
    .I1(net42),
    .S(_1540_),
    .Z(_0645_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1969_ (.I(_0645_),
    .Z(net148),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1970_ (.I0(\m_arbiter.wb0_o_dat[9] ),
    .I1(net43),
    .S(_1540_),
    .Z(_0646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1971_ (.I(_0646_),
    .Z(net149),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1972_ (.I0(\m_arbiter.wb0_o_dat[10] ),
    .I1(net29),
    .S(_1526_),
    .Z(_0647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1973_ (.I(_0647_),
    .Z(net135),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1974_ (.I0(\m_arbiter.wb0_o_dat[11] ),
    .I1(net30),
    .S(_1526_),
    .Z(_0648_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1975_ (.I(_0648_),
    .Z(net136),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1976_ (.I0(\m_arbiter.wb0_o_dat[12] ),
    .I1(net31),
    .S(_1540_),
    .Z(_0649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1977_ (.I(_0649_),
    .Z(net137),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1978_ (.I0(\m_arbiter.wb0_o_dat[13] ),
    .I1(net32),
    .S(_1540_),
    .Z(_0650_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1979_ (.I(_0650_),
    .Z(net138),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1980_ (.I0(\m_arbiter.wb0_o_dat[14] ),
    .I1(net33),
    .S(_1540_),
    .Z(_0651_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1981_ (.I(_0651_),
    .Z(net139),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1982_ (.I0(\m_arbiter.wb0_o_dat[15] ),
    .I1(net34),
    .S(_1540_),
    .Z(_0652_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1983_ (.I(_0652_),
    .Z(net140),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1984_ (.I0(clknet_leaf_50_user_clock2),
    .I1(\clk_div.res_clk ),
    .S(\clk_div.clock_sel_r ),
    .Z(_0653_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1985_ (.I(_0653_),
    .Z(net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1986_ (.A1(_1526_),
    .A2(net47),
    .ZN(_0654_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1987_ (.A1(_1524_),
    .A2(net499),
    .ZN(_0655_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1988_ (.A1(_0654_),
    .A2(_0655_),
    .ZN(_0656_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1989_ (.A1(_0591_),
    .A2(_0656_),
    .ZN(_0657_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1990_ (.I(_0657_),
    .ZN(_0658_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1991_ (.A1(_0457_),
    .A2(_0658_),
    .Z(_0659_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1992_ (.I(_0659_),
    .Z(net150),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1993_ (.I(_0542_),
    .Z(_0660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1994_ (.I(\wb_compressor.state[0] ),
    .ZN(_0661_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1995_ (.A1(_0660_),
    .A2(_0661_),
    .A3(_0575_),
    .ZN(_0001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1996_ (.A1(\wb_compressor.state[5] ),
    .A2(\wb_compressor.state[4] ),
    .ZN(_0662_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1997_ (.A1(_0543_),
    .A2(_0533_),
    .A3(_0540_),
    .A4(_0662_),
    .ZN(_0663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1998_ (.I(_0663_),
    .Z(_0000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1999_ (.A1(_1525_),
    .A2(_0596_),
    .ZN(net109),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2000_ (.A1(_1525_),
    .A2(_0590_),
    .ZN(net110),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2001_ (.A1(\wb_compressor.state[5] ),
    .A2(\wb_compressor.state[4] ),
    .B(_0533_),
    .ZN(_0664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2002_ (.A1(_0575_),
    .A2(_0662_),
    .ZN(_0665_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2003_ (.A1(\wb_compressor.state[6] ),
    .A2(\wb_compressor.state[2] ),
    .A3(_0555_),
    .ZN(_0666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2004_ (.A1(_0577_),
    .A2(_0664_),
    .A3(_0665_),
    .A4(_0666_),
    .Z(_0667_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2005_ (.I(_0667_),
    .Z(_0668_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2006_ (.A1(_0533_),
    .A2(_0662_),
    .ZN(_0669_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2007_ (.A1(_0540_),
    .A2(_0669_),
    .ZN(_0670_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2008_ (.A1(\wb_compressor.burst_cnt[0] ),
    .A2(_0668_),
    .ZN(_0671_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2009_ (.A1(_0668_),
    .A2(_0670_),
    .B(_0671_),
    .ZN(_0023_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2010_ (.A1(_0537_),
    .A2(_0536_),
    .A3(_0670_),
    .ZN(_0672_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2011_ (.I0(\wb_compressor.burst_cnt[1] ),
    .I1(_0672_),
    .S(_0668_),
    .Z(_0673_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2012_ (.I(_0673_),
    .Z(_0024_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2013_ (.A1(\wb_compressor.burst_cnt[2] ),
    .A2(_0536_),
    .A3(_0668_),
    .Z(_0674_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2014_ (.A1(_0536_),
    .A2(_0668_),
    .B(\wb_compressor.burst_cnt[2] ),
    .ZN(_0675_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2015_ (.A1(_0668_),
    .A2(_0670_),
    .B(_0674_),
    .C(_0675_),
    .ZN(_0025_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2016_ (.A1(\wb_compressor.wb_ack ),
    .A2(\wb_compressor.wb_err ),
    .ZN(_0676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2017_ (.I(_0676_),
    .Z(_0677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2018_ (.A1(_0521_),
    .A2(\wb_cross_clk.ack_xor_flag ),
    .Z(_0678_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2019_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[0] ),
    .A2(_0677_),
    .ZN(_0679_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2020_ (.A1(_0677_),
    .A2(_0678_),
    .B(_0679_),
    .ZN(_0026_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2021_ (.A1(\wb_compressor.wb_err ),
    .A2(\wb_cross_clk.err_xor_flag ),
    .ZN(_0680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2022_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[1] ),
    .A2(_0677_),
    .ZN(_0681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2023_ (.A1(_0677_),
    .A2(net245),
    .B(_0681_),
    .ZN(_0027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2024_ (.I0(\wb_compressor.wb_i_dat[0] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[2] ),
    .S(_0677_),
    .Z(_0682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2025_ (.I(_0682_),
    .Z(_0028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2026_ (.I0(\wb_compressor.wb_i_dat[1] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[3] ),
    .S(_0677_),
    .Z(_0683_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2027_ (.I(_0683_),
    .Z(_0029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2028_ (.I0(\wb_compressor.wb_i_dat[2] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[4] ),
    .S(_0677_),
    .Z(_0684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2029_ (.I(_0684_),
    .Z(_0030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2030_ (.I0(\wb_compressor.wb_i_dat[3] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[5] ),
    .S(_0677_),
    .Z(_0685_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2031_ (.I(_0685_),
    .Z(_0031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2032_ (.I0(\wb_compressor.wb_i_dat[4] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[6] ),
    .S(_0677_),
    .Z(_0686_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2033_ (.I(_0686_),
    .Z(_0032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2034_ (.I0(\wb_compressor.wb_i_dat[5] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[7] ),
    .S(_0677_),
    .Z(_0687_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2035_ (.I(_0687_),
    .Z(_0033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _2036_ (.I(_0676_),
    .Z(_0688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2037_ (.I0(\wb_compressor.wb_i_dat[6] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[8] ),
    .S(_0688_),
    .Z(_0689_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2038_ (.I(_0689_),
    .Z(_0034_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2039_ (.I0(\wb_compressor.wb_i_dat[7] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[9] ),
    .S(_0688_),
    .Z(_0690_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2040_ (.I(_0690_),
    .Z(_0035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2041_ (.I0(\wb_compressor.wb_i_dat[8] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[10] ),
    .S(_0688_),
    .Z(_0691_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2042_ (.I(_0691_),
    .Z(_0036_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2043_ (.I0(\wb_compressor.wb_i_dat[9] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[11] ),
    .S(_0688_),
    .Z(_0692_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2044_ (.I(_0692_),
    .Z(_0037_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2045_ (.I0(\wb_compressor.wb_i_dat[10] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[12] ),
    .S(_0688_),
    .Z(_0693_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2046_ (.I(_0693_),
    .Z(_0038_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2047_ (.I0(\wb_compressor.wb_i_dat[11] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[13] ),
    .S(_0688_),
    .Z(_0694_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2048_ (.I(_0694_),
    .Z(_0039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2049_ (.I0(\wb_compressor.wb_i_dat[12] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[14] ),
    .S(_0688_),
    .Z(_0695_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2050_ (.I(_0695_),
    .Z(_0040_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2051_ (.I0(\wb_compressor.wb_i_dat[13] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[15] ),
    .S(_0688_),
    .Z(_0696_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2052_ (.I(_0696_),
    .Z(_0041_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2053_ (.I0(\wb_compressor.wb_i_dat[14] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[16] ),
    .S(_0688_),
    .Z(_0697_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2054_ (.I(_0697_),
    .Z(_0042_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2055_ (.I0(\wb_compressor.wb_i_dat[15] ),
    .I1(\wb_cross_clk.s_m_sync.s_data_ff[17] ),
    .S(_0688_),
    .Z(_0698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2056_ (.I(_0698_),
    .Z(_0043_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _2057_ (.I(iram_wb_ack),
    .ZN(_0699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2058_ (.I(_0699_),
    .Z(_0700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2059_ (.A1(_0700_),
    .A2(_0457_),
    .A3(_0591_),
    .A4(_0596_),
    .Z(_0701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2060_ (.I(_0701_),
    .Z(_0044_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2061_ (.A1(_0700_),
    .A2(\iram_latched[0] ),
    .ZN(_0702_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2062_ (.I(iram_wb_ack),
    .Z(_0703_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2063_ (.A1(_0703_),
    .A2(net48),
    .ZN(_0704_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2064_ (.A1(_0702_),
    .A2(_0704_),
    .B(_0631_),
    .ZN(_0045_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2065_ (.A1(_0700_),
    .A2(\iram_latched[1] ),
    .ZN(_0705_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2066_ (.A1(_0703_),
    .A2(net55),
    .ZN(_0706_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2067_ (.A1(_0705_),
    .A2(_0706_),
    .B(_0631_),
    .ZN(_0046_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2068_ (.A1(_0700_),
    .A2(\iram_latched[2] ),
    .ZN(_0707_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2069_ (.A1(_0703_),
    .A2(net56),
    .ZN(_0708_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2070_ (.A1(_0707_),
    .A2(_0708_),
    .B(_0631_),
    .ZN(_0047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2071_ (.A1(_0700_),
    .A2(\iram_latched[3] ),
    .ZN(_0709_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2072_ (.A1(_0703_),
    .A2(net57),
    .ZN(_0710_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2073_ (.A1(_0709_),
    .A2(_0710_),
    .B(_0631_),
    .ZN(_0048_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2074_ (.A1(_0700_),
    .A2(\iram_latched[4] ),
    .ZN(_0711_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2075_ (.A1(_0703_),
    .A2(net58),
    .ZN(_0712_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2076_ (.A1(_0711_),
    .A2(_0712_),
    .B(_0631_),
    .ZN(_0049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2077_ (.A1(_0700_),
    .A2(\iram_latched[5] ),
    .ZN(_0713_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2078_ (.A1(_0703_),
    .A2(net59),
    .ZN(_0714_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2079_ (.A1(_0713_),
    .A2(_0714_),
    .B(_0631_),
    .ZN(_0050_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2080_ (.A1(_0700_),
    .A2(\iram_latched[6] ),
    .ZN(_0715_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2081_ (.A1(_0703_),
    .A2(net60),
    .ZN(_0716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2082_ (.A1(_0715_),
    .A2(_0716_),
    .B(_0631_),
    .ZN(_0051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2083_ (.A1(_0699_),
    .A2(\iram_latched[7] ),
    .ZN(_0717_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2084_ (.A1(_0703_),
    .A2(net61),
    .ZN(_0718_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2085_ (.A1(_0717_),
    .A2(_0718_),
    .B(_0631_),
    .ZN(_0052_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2086_ (.A1(_0699_),
    .A2(\iram_latched[8] ),
    .ZN(_0719_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2087_ (.A1(_0703_),
    .A2(net62),
    .ZN(_0720_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2088_ (.I(_0579_),
    .Z(_0721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2089_ (.A1(_0719_),
    .A2(_0720_),
    .B(_0721_),
    .ZN(_0053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2090_ (.A1(_0699_),
    .A2(\iram_latched[9] ),
    .ZN(_0722_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2091_ (.A1(iram_wb_ack),
    .A2(net63),
    .ZN(_0723_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2092_ (.A1(_0722_),
    .A2(_0723_),
    .B(_0721_),
    .ZN(_0054_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2093_ (.A1(_0699_),
    .A2(\iram_latched[10] ),
    .ZN(_0724_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2094_ (.A1(iram_wb_ack),
    .A2(net49),
    .ZN(_0725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2095_ (.A1(_0724_),
    .A2(_0725_),
    .B(_0721_),
    .ZN(_0055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2096_ (.A1(_0699_),
    .A2(\iram_latched[11] ),
    .ZN(_0726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2097_ (.A1(iram_wb_ack),
    .A2(net50),
    .ZN(_0727_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2098_ (.A1(_0726_),
    .A2(_0727_),
    .B(_0721_),
    .ZN(_0056_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2099_ (.A1(_0699_),
    .A2(\iram_latched[12] ),
    .ZN(_0728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2100_ (.A1(iram_wb_ack),
    .A2(net51),
    .ZN(_0729_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2101_ (.A1(_0728_),
    .A2(_0729_),
    .B(_0721_),
    .ZN(_0057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2102_ (.A1(_0699_),
    .A2(\iram_latched[13] ),
    .ZN(_0730_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2103_ (.A1(iram_wb_ack),
    .A2(net52),
    .ZN(_0731_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2104_ (.A1(_0730_),
    .A2(_0731_),
    .B(_0721_),
    .ZN(_0058_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2105_ (.A1(_0699_),
    .A2(\iram_latched[14] ),
    .ZN(_0732_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2106_ (.A1(iram_wb_ack),
    .A2(net53),
    .ZN(_0733_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2107_ (.A1(_0732_),
    .A2(_0733_),
    .B(_0721_),
    .ZN(_0059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2108_ (.A1(\iram_latched[15] ),
    .A2(_0700_),
    .ZN(_0734_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2109_ (.A1(net54),
    .A2(_0703_),
    .ZN(_0735_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2110_ (.A1(_0734_),
    .A2(_0735_),
    .B(_0721_),
    .ZN(_0060_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2111_ (.A1(_0700_),
    .A2(_0631_),
    .ZN(_0061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2112_ (.I(\clk_div.curr_div[2] ),
    .ZN(_0736_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2113_ (.I(\clk_div.curr_div[0] ),
    .Z(_0737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2114_ (.I0(\clk_div.cnt[8] ),
    .I1(\clk_div.cnt[9] ),
    .I2(\clk_div.cnt[10] ),
    .I3(\clk_div.cnt[11] ),
    .S0(_0737_),
    .S1(\clk_div.curr_div[1] ),
    .Z(_0738_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2115_ (.A1(_0736_),
    .A2(_0738_),
    .ZN(_0739_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _2116_ (.I0(\clk_div.cnt[12] ),
    .I1(\clk_div.cnt[13] ),
    .I2(\clk_div.cnt[14] ),
    .I3(\clk_div.cnt[15] ),
    .S0(_0737_),
    .S1(\clk_div.curr_div[1] ),
    .Z(_0740_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2117_ (.I(\clk_div.curr_div[3] ),
    .ZN(_0741_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2118_ (.A1(\clk_div.curr_div[2] ),
    .A2(_0740_),
    .B(_0741_),
    .ZN(_0742_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2119_ (.I0(\clk_div.cnt[4] ),
    .I1(\clk_div.cnt[5] ),
    .I2(\clk_div.cnt[6] ),
    .I3(\clk_div.cnt[7] ),
    .S0(_0737_),
    .S1(\clk_div.curr_div[1] ),
    .Z(_0743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2120_ (.A1(\clk_div.curr_div[2] ),
    .A2(_0743_),
    .B(\clk_div.curr_div[3] ),
    .ZN(_0744_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2121_ (.I0(\clk_div.cnt[0] ),
    .I1(\clk_div.cnt[1] ),
    .I2(\clk_div.cnt[2] ),
    .I3(\clk_div.cnt[3] ),
    .S0(_0737_),
    .S1(\clk_div.curr_div[1] ),
    .Z(_0745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2122_ (.A1(_0736_),
    .A2(_0745_),
    .ZN(_0746_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2123_ (.A1(_0739_),
    .A2(_0742_),
    .B1(_0744_),
    .B2(_0746_),
    .ZN(_0747_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2124_ (.A1(\clk_div.res_clk ),
    .A2(net244),
    .Z(_0748_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2125_ (.I(_0748_),
    .Z(_0062_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2126_ (.A1(_1570_),
    .A2(_0394_),
    .A3(net255),
    .A4(_0397_),
    .ZN(_0749_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2127_ (.A1(_0469_),
    .A2(_0407_),
    .A3(_0409_),
    .A4(_0749_),
    .ZN(_0750_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2128_ (.A1(_0750_),
    .A2(_0525_),
    .A3(_0656_),
    .ZN(_0751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2129_ (.A1(\clk_div.next_div_buff[0] ),
    .A2(_0751_),
    .ZN(_0752_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2130_ (.A1(_1552_),
    .A2(_0751_),
    .B(_0752_),
    .ZN(_0063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2131_ (.A1(\clk_div.next_div_buff[1] ),
    .A2(_0751_),
    .ZN(_0753_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2132_ (.A1(_1548_),
    .A2(_0751_),
    .B(_0753_),
    .ZN(_0064_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2133_ (.A1(\clk_div.next_div_buff[2] ),
    .A2(_0751_),
    .ZN(_0754_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2134_ (.A1(_1544_),
    .A2(_0751_),
    .B(_0754_),
    .ZN(_0065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2135_ (.A1(\clk_div.next_div_buff[3] ),
    .A2(_0751_),
    .ZN(_0755_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2136_ (.A1(_1539_),
    .A2(_0751_),
    .B(_0755_),
    .ZN(_0066_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2137_ (.I(_0747_),
    .ZN(_0756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2138_ (.A1(\clk_div.next_div_val ),
    .A2(_0756_),
    .ZN(_0757_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2139_ (.A1(_0751_),
    .A2(_0757_),
    .B(_0721_),
    .ZN(_0067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2140_ (.I(\clk_div.next_div_buff[0] ),
    .ZN(_0758_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2141_ (.A1(\clk_div.next_div_val ),
    .A2(_0747_),
    .ZN(_0759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2142_ (.A1(_0737_),
    .A2(_0759_),
    .ZN(_0760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2143_ (.I(_0622_),
    .Z(_0761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2144_ (.A1(_0758_),
    .A2(_0759_),
    .B(_0760_),
    .C(_0761_),
    .ZN(_0068_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2145_ (.I(\clk_div.curr_div[1] ),
    .ZN(_0762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2146_ (.I(_0622_),
    .Z(_0763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2147_ (.A1(\clk_div.next_div_buff[1] ),
    .A2(_0759_),
    .B(_0763_),
    .ZN(_0764_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2148_ (.A1(_0762_),
    .A2(_0759_),
    .B(_0764_),
    .ZN(_0069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2149_ (.I(\clk_div.next_div_buff[2] ),
    .ZN(_0765_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2150_ (.A1(\clk_div.curr_div[2] ),
    .A2(_0759_),
    .ZN(_0766_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2151_ (.A1(_0765_),
    .A2(_0759_),
    .B(_0766_),
    .C(_0761_),
    .ZN(_0070_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2152_ (.A1(\clk_div.next_div_buff[3] ),
    .A2(_0759_),
    .B(_0763_),
    .ZN(_0767_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2153_ (.A1(_0741_),
    .A2(_0759_),
    .B(_0767_),
    .ZN(_0071_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2154_ (.I(\wb_cross_clk.m_s_sync.d_data[0] ),
    .ZN(_0768_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2155_ (.I(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[1] ),
    .ZN(_0769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2156_ (.A1(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[2] ),
    .A2(_0769_),
    .Z(_0770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2157_ (.I(_0770_),
    .Z(_0771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2158_ (.I(_0770_),
    .Z(_0772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2159_ (.A1(net482),
    .A2(_0772_),
    .ZN(_0773_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2160_ (.I(_0542_),
    .Z(_0774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2161_ (.A1(_0768_),
    .A2(_0771_),
    .B(_0773_),
    .C(_0774_),
    .ZN(_0072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2162_ (.A1(\wb_cross_clk.m_s_sync.d_data[1] ),
    .A2(_0771_),
    .ZN(_0775_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _2163_ (.A1(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[2] ),
    .A2(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[1] ),
    .Z(_0776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2164_ (.I(_0776_),
    .Z(_0777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2165_ (.A1(net412),
    .A2(_0777_),
    .ZN(_0778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2166_ (.A1(_0775_),
    .A2(net413),
    .B(_0544_),
    .ZN(_0073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2167_ (.I(net480),
    .ZN(_0779_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2168_ (.A1(\wb_cross_clk.m_s_sync.d_data[2] ),
    .A2(_0776_),
    .ZN(_0780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2169_ (.A1(net481),
    .A2(_0777_),
    .B(_0780_),
    .C(_0774_),
    .ZN(_0074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2170_ (.A1(\wb_cross_clk.m_s_sync.d_data[3] ),
    .A2(_0771_),
    .ZN(_0781_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2171_ (.A1(net426),
    .A2(_0777_),
    .ZN(_0782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2172_ (.A1(_0781_),
    .A2(net427),
    .B(_0544_),
    .ZN(_0075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2173_ (.I(_0770_),
    .Z(_0783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2174_ (.A1(\wb_cross_clk.m_s_sync.d_data[4] ),
    .A2(_0783_),
    .ZN(_0784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2175_ (.A1(net442),
    .A2(_0777_),
    .ZN(_0785_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2176_ (.A1(_0784_),
    .A2(net443),
    .B(_0544_),
    .ZN(_0076_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2177_ (.A1(\wb_cross_clk.m_s_sync.d_data[5] ),
    .A2(_0783_),
    .ZN(_0786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2178_ (.A1(net444),
    .A2(_0777_),
    .ZN(_0787_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2179_ (.A1(_0786_),
    .A2(net445),
    .B(_0544_),
    .ZN(_0077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2180_ (.A1(\wb_cross_clk.m_s_sync.d_data[6] ),
    .A2(_0783_),
    .ZN(_0788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2181_ (.A1(net432),
    .A2(_0777_),
    .ZN(_0789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2182_ (.A1(_0788_),
    .A2(net433),
    .B(_0544_),
    .ZN(_0078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2183_ (.A1(\wb_cross_clk.m_s_sync.d_data[7] ),
    .A2(_0783_),
    .ZN(_0790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2184_ (.A1(net416),
    .A2(_0777_),
    .ZN(_0791_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2185_ (.A1(_0790_),
    .A2(net417),
    .B(_0544_),
    .ZN(_0079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2186_ (.A1(\wb_cross_clk.m_s_sync.d_data[8] ),
    .A2(_0783_),
    .ZN(_0792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2187_ (.A1(net418),
    .A2(_0777_),
    .ZN(_0793_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2188_ (.I(_0543_),
    .Z(_0794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2189_ (.A1(_0792_),
    .A2(net419),
    .B(_0794_),
    .ZN(_0080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2190_ (.A1(\wb_cross_clk.m_s_sync.d_data[9] ),
    .A2(_0783_),
    .ZN(_0795_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2191_ (.A1(net404),
    .A2(_0777_),
    .ZN(_0796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2192_ (.A1(_0795_),
    .A2(net405),
    .B(_0794_),
    .ZN(_0081_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2193_ (.A1(\wb_cross_clk.m_s_sync.d_data[10] ),
    .A2(_0783_),
    .ZN(_0797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2194_ (.A1(net428),
    .A2(_0777_),
    .ZN(_0798_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2195_ (.A1(_0797_),
    .A2(net429),
    .B(_0794_),
    .ZN(_0082_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2196_ (.A1(\wb_cross_clk.m_s_sync.d_data[11] ),
    .A2(_0783_),
    .ZN(_0799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2197_ (.I(_0776_),
    .Z(_0800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2198_ (.A1(net414),
    .A2(_0800_),
    .ZN(_0801_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2199_ (.A1(_0799_),
    .A2(net415),
    .B(_0794_),
    .ZN(_0083_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2200_ (.A1(\wb_cross_clk.m_s_sync.d_data[12] ),
    .A2(_0783_),
    .ZN(_0802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2201_ (.A1(net452),
    .A2(_0800_),
    .ZN(_0803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2202_ (.A1(_0802_),
    .A2(net453),
    .B(_0794_),
    .ZN(_0084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2203_ (.A1(\wb_cross_clk.m_s_sync.d_data[13] ),
    .A2(_0783_),
    .ZN(_0804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2204_ (.A1(net450),
    .A2(_0800_),
    .ZN(_0805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2205_ (.A1(_0804_),
    .A2(net451),
    .B(_0794_),
    .ZN(_0085_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2206_ (.I(_0770_),
    .Z(_0806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2207_ (.A1(\wb_cross_clk.m_s_sync.d_data[14] ),
    .A2(_0806_),
    .ZN(_0807_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2208_ (.A1(net408),
    .A2(_0800_),
    .ZN(_0808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2209_ (.A1(_0807_),
    .A2(net409),
    .B(_0794_),
    .ZN(_0086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2210_ (.A1(\wb_cross_clk.m_s_sync.d_data[15] ),
    .A2(_0806_),
    .ZN(_0809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2211_ (.A1(net434),
    .A2(_0800_),
    .ZN(_0810_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2212_ (.A1(_0809_),
    .A2(net435),
    .B(_0794_),
    .ZN(_0087_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2213_ (.A1(\wb_cross_clk.m_s_sync.d_data[16] ),
    .A2(_0806_),
    .ZN(_0811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2214_ (.A1(net474),
    .A2(_0800_),
    .ZN(_0812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2215_ (.A1(_0811_),
    .A2(net475),
    .B(_0794_),
    .ZN(_0088_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2216_ (.A1(\wb_cross_clk.m_s_sync.d_data[17] ),
    .A2(_0806_),
    .ZN(_0813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2217_ (.A1(net454),
    .A2(_0800_),
    .ZN(_0814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2218_ (.A1(_0813_),
    .A2(net455),
    .B(_0794_),
    .ZN(_0089_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2219_ (.A1(\wb_cross_clk.m_s_sync.d_data[18] ),
    .A2(_0806_),
    .ZN(_0815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2220_ (.A1(net424),
    .A2(_0800_),
    .ZN(_0816_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2221_ (.I(_0543_),
    .Z(_0817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2222_ (.A1(_0815_),
    .A2(net425),
    .B(_0817_),
    .ZN(_0090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2223_ (.I(\wb_cross_clk.m_s_sync.d_data[19] ),
    .ZN(_0818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2224_ (.A1(net483),
    .A2(_0772_),
    .ZN(_0819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2225_ (.A1(_0818_),
    .A2(_0771_),
    .B(_0819_),
    .C(_0774_),
    .ZN(_0091_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2226_ (.I(\wb_cross_clk.m_s_sync.d_data[20] ),
    .ZN(_0820_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2227_ (.A1(net484),
    .A2(_0772_),
    .ZN(_0821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2228_ (.A1(_0820_),
    .A2(_0771_),
    .B(_0821_),
    .C(_0774_),
    .ZN(_0092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2229_ (.I(\wb_cross_clk.m_s_sync.d_data[21] ),
    .ZN(_0822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2230_ (.A1(net485),
    .A2(_0772_),
    .ZN(_0823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2231_ (.A1(_0822_),
    .A2(_0771_),
    .B(_0823_),
    .C(_0660_),
    .ZN(_0093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2232_ (.A1(\wb_cross_clk.m_s_sync.d_data[22] ),
    .A2(_0806_),
    .ZN(_0824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2233_ (.A1(net422),
    .A2(_0800_),
    .ZN(_0825_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2234_ (.A1(_0824_),
    .A2(net423),
    .B(_0817_),
    .ZN(_0094_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2235_ (.A1(\wb_cross_clk.m_s_sync.d_data[23] ),
    .A2(_0806_),
    .ZN(_0826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2236_ (.A1(net430),
    .A2(_0800_),
    .ZN(_0827_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2237_ (.A1(_0826_),
    .A2(net431),
    .B(_0817_),
    .ZN(_0095_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2238_ (.A1(\wb_cross_clk.m_s_sync.d_data[24] ),
    .A2(_0806_),
    .ZN(_0828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2239_ (.I(_0776_),
    .Z(_0829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2240_ (.A1(net440),
    .A2(_0829_),
    .ZN(_0830_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2241_ (.A1(_0828_),
    .A2(net441),
    .B(_0817_),
    .ZN(_0096_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2242_ (.A1(\wb_cross_clk.m_s_sync.d_data[25] ),
    .A2(_0806_),
    .ZN(_0831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2243_ (.A1(net410),
    .A2(_0829_),
    .ZN(_0832_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2244_ (.A1(_0831_),
    .A2(net411),
    .B(_0817_),
    .ZN(_0097_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2245_ (.A1(\wb_cross_clk.m_s_sync.d_data[26] ),
    .A2(_0806_),
    .ZN(_0833_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2246_ (.A1(net398),
    .A2(_0829_),
    .ZN(_0834_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2247_ (.A1(_0833_),
    .A2(net399),
    .B(_0817_),
    .ZN(_0098_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2248_ (.I(_0770_),
    .Z(_0835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2249_ (.A1(\wb_cross_clk.m_s_sync.d_data[27] ),
    .A2(_0835_),
    .ZN(_0836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2250_ (.A1(net462),
    .A2(_0829_),
    .ZN(_0837_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2251_ (.A1(_0836_),
    .A2(net463),
    .B(_0817_),
    .ZN(_0099_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2252_ (.A1(\wb_cross_clk.m_s_sync.d_data[28] ),
    .A2(_0835_),
    .ZN(_0838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2253_ (.A1(net420),
    .A2(_0829_),
    .ZN(_0839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2254_ (.A1(_0838_),
    .A2(net421),
    .B(_0817_),
    .ZN(_0100_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2255_ (.A1(\wb_cross_clk.m_s_sync.d_data[29] ),
    .A2(_0835_),
    .ZN(_0840_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2256_ (.A1(net472),
    .A2(_0829_),
    .ZN(_0841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2257_ (.A1(_0840_),
    .A2(net473),
    .B(_0817_),
    .ZN(_0101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2258_ (.A1(\wb_cross_clk.m_s_sync.d_data[30] ),
    .A2(_0835_),
    .ZN(_0842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2259_ (.A1(net396),
    .A2(_0829_),
    .ZN(_0843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2260_ (.A1(_0842_),
    .A2(net397),
    .B(_0817_),
    .ZN(_0102_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2261_ (.A1(\wb_cross_clk.m_s_sync.d_data[31] ),
    .A2(_0835_),
    .ZN(_0844_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2262_ (.A1(net456),
    .A2(_0829_),
    .ZN(_0845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2263_ (.I(_0543_),
    .Z(_0846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2264_ (.A1(_0844_),
    .A2(net457),
    .B(_0846_),
    .ZN(_0103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2265_ (.A1(\wb_cross_clk.m_s_sync.d_data[32] ),
    .A2(_0835_),
    .ZN(_0847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2266_ (.A1(net464),
    .A2(_0829_),
    .ZN(_0848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2267_ (.A1(_0847_),
    .A2(net465),
    .B(_0846_),
    .ZN(_0104_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2268_ (.A1(\wb_cross_clk.m_s_sync.d_data[33] ),
    .A2(_0835_),
    .ZN(_0849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2269_ (.A1(net448),
    .A2(_0829_),
    .ZN(_0850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2270_ (.A1(_0849_),
    .A2(net449),
    .B(_0846_),
    .ZN(_0105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2271_ (.A1(\wb_cross_clk.m_s_sync.d_data[34] ),
    .A2(_0835_),
    .ZN(_0851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2272_ (.I(_0776_),
    .Z(_0852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2273_ (.A1(net436),
    .A2(_0852_),
    .ZN(_0853_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2274_ (.A1(_0851_),
    .A2(net437),
    .B(_0846_),
    .ZN(_0106_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2275_ (.A1(\wb_cross_clk.m_s_sync.d_data[35] ),
    .A2(_0835_),
    .ZN(_0854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2276_ (.A1(net438),
    .A2(_0852_),
    .ZN(_0855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2277_ (.A1(_0854_),
    .A2(net439),
    .B(_0846_),
    .ZN(_0107_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2278_ (.A1(\wb_cross_clk.m_s_sync.d_data[36] ),
    .A2(_0835_),
    .ZN(_0856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2279_ (.A1(net446),
    .A2(_0852_),
    .ZN(_0857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2280_ (.A1(_0856_),
    .A2(net447),
    .B(_0846_),
    .ZN(_0108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2281_ (.A1(\wb_cross_clk.m_s_sync.d_data[37] ),
    .A2(_0772_),
    .ZN(_0858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2282_ (.A1(net476),
    .A2(_0852_),
    .ZN(_0859_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2283_ (.A1(_0858_),
    .A2(net477),
    .B(_0846_),
    .ZN(_0109_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2284_ (.A1(net466),
    .A2(_0852_),
    .ZN(_0860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2285_ (.A1(\wb_cross_clk.m_s_sync.d_data[38] ),
    .A2(_0771_),
    .ZN(_0861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2286_ (.A1(net467),
    .A2(_0861_),
    .B(_0846_),
    .ZN(_0110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2287_ (.A1(net406),
    .A2(_0776_),
    .ZN(_0862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2288_ (.A1(\wb_cross_clk.m_s_sync.d_data[39] ),
    .A2(_0771_),
    .ZN(_0863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2289_ (.A1(net407),
    .A2(_0863_),
    .B(_0846_),
    .ZN(_0111_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2290_ (.A1(\wb_cross_clk.m_s_sync.d_data[40] ),
    .A2(_0772_),
    .ZN(_0864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2291_ (.A1(net402),
    .A2(_0852_),
    .ZN(_0865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2292_ (.A1(_0864_),
    .A2(net403),
    .B(_0846_),
    .ZN(_0112_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2293_ (.A1(net394),
    .A2(_0776_),
    .ZN(_0866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2294_ (.A1(\wb_cross_clk.m_s_sync.d_data[41] ),
    .A2(_0771_),
    .ZN(_0867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2295_ (.A1(net395),
    .A2(_0867_),
    .B(_0549_),
    .ZN(_0113_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2296_ (.A1(net460),
    .A2(_0776_),
    .ZN(_0868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2297_ (.A1(\wb_cross_clk.m_s_sync.d_data[42] ),
    .A2(_0771_),
    .ZN(_0869_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2298_ (.A1(net461),
    .A2(_0869_),
    .B(_0549_),
    .ZN(_0114_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2299_ (.A1(\wb_cross_clk.m_s_sync.d_data[43] ),
    .A2(_0772_),
    .ZN(_0870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2300_ (.A1(net478),
    .A2(_0852_),
    .ZN(_0871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2301_ (.A1(_0870_),
    .A2(net479),
    .B(_0549_),
    .ZN(_0115_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2302_ (.A1(\wb_cross_clk.m_s_sync.d_data[44] ),
    .A2(_0772_),
    .ZN(_0872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2303_ (.A1(net468),
    .A2(_0852_),
    .ZN(_0873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2304_ (.A1(_0872_),
    .A2(net469),
    .B(_0549_),
    .ZN(_0116_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2305_ (.A1(\wb_cross_clk.m_s_sync.d_data[45] ),
    .A2(_0772_),
    .ZN(_0874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2306_ (.A1(net470),
    .A2(_0852_),
    .ZN(_0875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2307_ (.A1(_0874_),
    .A2(net471),
    .B(_0549_),
    .ZN(_0117_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2308_ (.A1(\wb_cross_clk.m_s_sync.d_data[46] ),
    .A2(_0772_),
    .ZN(_0876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2309_ (.A1(net458),
    .A2(_0852_),
    .ZN(_0877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2310_ (.A1(_0876_),
    .A2(net459),
    .B(_0549_),
    .ZN(_0118_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2311_ (.A1(net262),
    .A2(net260),
    .Z(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2312_ (.A1(_0634_),
    .A2(_0878_),
    .ZN(_0119_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2313_ (.I(net400),
    .ZN(_0879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2314_ (.A1(_1540_),
    .A2(\m_arbiter.i_wb0_cyc ),
    .B(_0412_),
    .C(_0526_),
    .ZN(_0880_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2315_ (.I(\wb_cross_clk.prev_stb ),
    .ZN(_0881_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2316_ (.A1(\wb_cross_clk.m_burst_cnt[3] ),
    .A2(\wb_cross_clk.m_burst_cnt[2] ),
    .A3(\wb_cross_clk.m_burst_cnt[1] ),
    .A4(\wb_cross_clk.m_burst_cnt[0] ),
    .ZN(_0882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2317_ (.A1(_0881_),
    .A2(\wb_cross_clk.prev_ack ),
    .B(_0882_),
    .ZN(_0883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2318_ (.A1(_0394_),
    .A2(_0395_),
    .B(_0880_),
    .C(_0883_),
    .ZN(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2319_ (.I(net210),
    .Z(_0885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2320_ (.A1(_0879_),
    .A2(_0885_),
    .Z(_0886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2321_ (.A1(_0634_),
    .A2(_0886_),
    .ZN(_0120_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2322_ (.A1(net401),
    .A2(_0544_),
    .ZN(_0121_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2323_ (.I(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[0] ),
    .ZN(_0887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2324_ (.A1(_0553_),
    .A2(_0887_),
    .ZN(_0122_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2325_ (.A1(_0553_),
    .A2(_0769_),
    .ZN(_0123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _2326_ (.A1(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[2] ),
    .A2(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[1] ),
    .ZN(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2327_ (.I(_0888_),
    .Z(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2328_ (.A1(\wb_cross_clk.msy_xor_ack ),
    .A2(_0889_),
    .ZN(_0890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _2329_ (.A1(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[2] ),
    .A2(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[1] ),
    .Z(_0891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2330_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[0] ),
    .A2(_0891_),
    .ZN(_0892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2331_ (.A1(_0890_),
    .A2(_0892_),
    .B(_0721_),
    .ZN(_0124_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2332_ (.A1(\wb_cross_clk.msy_xor_err ),
    .A2(_0889_),
    .ZN(_0893_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2333_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[1] ),
    .A2(_0891_),
    .ZN(_0894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2334_ (.I(_0579_),
    .Z(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2335_ (.A1(_0893_),
    .A2(_0894_),
    .B(_0895_),
    .ZN(_0125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2336_ (.I(_0888_),
    .Z(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2337_ (.A1(\wb_cross_clk.m_wb_i_dat[0] ),
    .A2(_0896_),
    .ZN(_0897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2338_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[2] ),
    .A2(_0891_),
    .ZN(_0898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2339_ (.A1(_0897_),
    .A2(_0898_),
    .B(_0895_),
    .ZN(_0126_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2340_ (.A1(\wb_cross_clk.m_wb_i_dat[1] ),
    .A2(_0896_),
    .ZN(_0899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2341_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[3] ),
    .A2(_0891_),
    .ZN(_0900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2342_ (.A1(_0899_),
    .A2(_0900_),
    .B(_0895_),
    .ZN(_0127_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2343_ (.A1(\wb_cross_clk.m_wb_i_dat[2] ),
    .A2(_0896_),
    .ZN(_0901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2344_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[4] ),
    .A2(_0891_),
    .ZN(_0902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2345_ (.A1(_0901_),
    .A2(_0902_),
    .B(_0895_),
    .ZN(_0128_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2346_ (.A1(\wb_cross_clk.m_wb_i_dat[3] ),
    .A2(_0896_),
    .ZN(_0903_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2347_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[5] ),
    .A2(_0891_),
    .ZN(_0904_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2348_ (.A1(_0903_),
    .A2(_0904_),
    .B(_0895_),
    .ZN(_0129_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2349_ (.A1(\wb_cross_clk.m_wb_i_dat[4] ),
    .A2(_0896_),
    .ZN(_0905_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2350_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[6] ),
    .A2(_0891_),
    .ZN(_0906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2351_ (.A1(_0905_),
    .A2(_0906_),
    .B(_0895_),
    .ZN(_0130_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2352_ (.A1(\wb_cross_clk.m_wb_i_dat[5] ),
    .A2(_0896_),
    .ZN(_0907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2353_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[7] ),
    .A2(_0891_),
    .ZN(_0908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2354_ (.A1(_0907_),
    .A2(_0908_),
    .B(_0895_),
    .ZN(_0131_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2355_ (.A1(\wb_cross_clk.m_wb_i_dat[6] ),
    .A2(_0896_),
    .ZN(_0909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2356_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[8] ),
    .A2(_0891_),
    .ZN(_0910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2357_ (.A1(_0909_),
    .A2(_0910_),
    .B(_0895_),
    .ZN(_0132_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2358_ (.A1(\wb_cross_clk.m_wb_i_dat[7] ),
    .A2(_0896_),
    .ZN(_0911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2359_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[9] ),
    .A2(_0891_),
    .ZN(_0912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2360_ (.A1(_0911_),
    .A2(_0912_),
    .B(_0895_),
    .ZN(_0133_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2361_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[10] ),
    .A2(_0896_),
    .ZN(_0913_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2362_ (.A1(_0453_),
    .A2(_0889_),
    .B(_0913_),
    .C(_0580_),
    .ZN(_0134_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2363_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[11] ),
    .A2(_0896_),
    .ZN(_0914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2364_ (.A1(_0449_),
    .A2(_0889_),
    .B(_0914_),
    .C(_0580_),
    .ZN(_0135_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2365_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[12] ),
    .A2(_0888_),
    .ZN(_0915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2366_ (.A1(_0445_),
    .A2(_0889_),
    .B(_0915_),
    .C(_0580_),
    .ZN(_0136_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2367_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[13] ),
    .A2(_0888_),
    .ZN(_0916_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2368_ (.I(_0579_),
    .Z(_0917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2369_ (.A1(_0441_),
    .A2(_0889_),
    .B(_0916_),
    .C(_0917_),
    .ZN(_0137_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2370_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[14] ),
    .A2(_0888_),
    .ZN(_0918_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2371_ (.A1(_0437_),
    .A2(_0889_),
    .B(_0918_),
    .C(_0917_),
    .ZN(_0138_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2372_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[15] ),
    .A2(_0888_),
    .ZN(_0919_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2373_ (.A1(_0433_),
    .A2(_0889_),
    .B(_0919_),
    .C(_0917_),
    .ZN(_0139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2374_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[16] ),
    .A2(_0888_),
    .ZN(_0920_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2375_ (.A1(_0429_),
    .A2(_0889_),
    .B(_0920_),
    .C(_0917_),
    .ZN(_0140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2376_ (.A1(\wb_cross_clk.s_m_sync.s_data_ff[17] ),
    .A2(_0888_),
    .ZN(_0921_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2377_ (.A1(_0414_),
    .A2(_0889_),
    .B(_0921_),
    .C(_0917_),
    .ZN(_0141_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2378_ (.I(\wb_cross_clk.m_new_req_flag ),
    .ZN(_0922_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _2379_ (.I(net209),
    .Z(_0923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2380_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[0] ),
    .I1(_0922_),
    .S(_0923_),
    .Z(_0924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2381_ (.I(_0924_),
    .Z(_0142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2382_ (.I(_0885_),
    .Z(_0925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2383_ (.A1(_1540_),
    .A2(net2),
    .ZN(_0926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2384_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[1] ),
    .A2(_0925_),
    .ZN(_0927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2385_ (.A1(_0925_),
    .A2(_0926_),
    .B(_0927_),
    .ZN(_0143_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2386_ (.A1(_1527_),
    .A2(net1),
    .A3(net210),
    .ZN(_0928_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2387_ (.A1(_0779_),
    .A2(_0925_),
    .B(_0928_),
    .ZN(_0144_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2388_ (.A1(_1525_),
    .A2(net44),
    .Z(_0929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2389_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[3] ),
    .I1(_0929_),
    .S(_0923_),
    .Z(_0930_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2390_ (.I(_0930_),
    .Z(_0145_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2391_ (.A1(_1525_),
    .A2(net45),
    .Z(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2392_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[4] ),
    .I1(_0931_),
    .S(_0923_),
    .Z(_0932_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2393_ (.I(_0932_),
    .Z(_0146_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2394_ (.A1(_0654_),
    .A2(_0655_),
    .Z(_0933_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2395_ (.I(_0885_),
    .Z(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2396_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[5] ),
    .A2(_0925_),
    .ZN(_0935_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2397_ (.A1(_0933_),
    .A2(_0934_),
    .B(_0935_),
    .ZN(_0147_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2398_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[6] ),
    .A2(_0925_),
    .ZN(_0936_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2399_ (.A1(_1552_),
    .A2(_0934_),
    .B(_0936_),
    .ZN(_0148_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2400_ (.I(_0885_),
    .Z(_0937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2401_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[7] ),
    .A2(_0937_),
    .ZN(_0938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2402_ (.A1(_1548_),
    .A2(_0934_),
    .B(_0938_),
    .ZN(_0149_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2403_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[8] ),
    .A2(_0937_),
    .ZN(_0939_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2404_ (.A1(_1544_),
    .A2(_0934_),
    .B(_0939_),
    .ZN(_0150_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2405_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[9] ),
    .A2(_0937_),
    .ZN(_0940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2406_ (.A1(_1539_),
    .A2(_0934_),
    .B(_0940_),
    .ZN(_0151_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2407_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[10] ),
    .A2(_0937_),
    .ZN(_0941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2408_ (.A1(net234),
    .A2(_0934_),
    .B(_0941_),
    .ZN(_0152_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2409_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[11] ),
    .A2(_0937_),
    .ZN(_0942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2410_ (.A1(net235),
    .A2(_0934_),
    .B(_0942_),
    .ZN(_0153_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2411_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[12] ),
    .A2(_0937_),
    .ZN(_0943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2412_ (.A1(net236),
    .A2(_0934_),
    .B(_0943_),
    .ZN(_0154_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2413_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[13] ),
    .A2(_0937_),
    .ZN(_0944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2414_ (.A1(net237),
    .A2(_0934_),
    .B(_0944_),
    .ZN(_0155_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2415_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[14] ),
    .I1(net148),
    .S(_0923_),
    .Z(_0945_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2416_ (.I(_0945_),
    .Z(_0156_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2417_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[15] ),
    .I1(net149),
    .S(_0923_),
    .Z(_0946_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2418_ (.I(_0946_),
    .Z(_0157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2419_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[16] ),
    .I1(net135),
    .S(_0923_),
    .Z(_0947_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2420_ (.I(_0947_),
    .Z(_0158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2421_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[17] ),
    .I1(net136),
    .S(_0923_),
    .Z(_0948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2422_ (.I(_0948_),
    .Z(_0159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _2423_ (.I(net211),
    .Z(_0949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2424_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[18] ),
    .I1(net137),
    .S(_0949_),
    .Z(_0950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2425_ (.I(_0950_),
    .Z(_0160_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2426_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[19] ),
    .I1(net138),
    .S(_0949_),
    .Z(_0951_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2427_ (.I(_0951_),
    .Z(_0161_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2428_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[20] ),
    .I1(net139),
    .S(_0949_),
    .Z(_0952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2429_ (.I(_0952_),
    .Z(_0162_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2430_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[21] ),
    .I1(net140),
    .S(_0949_),
    .Z(_0953_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2431_ (.I(_0953_),
    .Z(_0163_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2432_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[22] ),
    .A2(_0937_),
    .ZN(_0954_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2433_ (.A1(_0463_),
    .A2(_0934_),
    .B(_0954_),
    .ZN(_0164_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2434_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[23] ),
    .A2(_0937_),
    .ZN(_0955_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2435_ (.A1(_0408_),
    .A2(_0925_),
    .B(_0955_),
    .ZN(_0165_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2436_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[24] ),
    .I1(net129),
    .S(_0949_),
    .Z(_0956_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2437_ (.I(_0956_),
    .Z(_0166_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2438_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[25] ),
    .I1(net130),
    .S(_0949_),
    .Z(_0957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2439_ (.I(_0957_),
    .Z(_0167_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2440_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[26] ),
    .A2(_0937_),
    .ZN(_0958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2441_ (.A1(_1593_),
    .A2(_0925_),
    .B(_0958_),
    .ZN(_0168_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2442_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[27] ),
    .A2(_0923_),
    .ZN(_0959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2443_ (.A1(_0406_),
    .A2(_0925_),
    .B(_0959_),
    .ZN(_0169_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2444_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[28] ),
    .I1(_1564_),
    .S(_0949_),
    .Z(_0960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2445_ (.I(_0960_),
    .Z(_0170_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2446_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[29] ),
    .I1(_1563_),
    .S(_0949_),
    .Z(_0961_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2447_ (.I(_0961_),
    .Z(_0171_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2448_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[30] ),
    .I1(_0396_),
    .S(_0949_),
    .Z(_0962_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2449_ (.I(_0962_),
    .Z(_0172_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2450_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[31] ),
    .I1(_1558_),
    .S(_0949_),
    .Z(_0963_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2451_ (.I(_0963_),
    .Z(_0173_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _2452_ (.I(net211),
    .Z(_0964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2453_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[32] ),
    .I1(_1582_),
    .S(_0964_),
    .Z(_0965_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2454_ (.I(_0965_),
    .Z(_0174_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2455_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[33] ),
    .I1(_1581_),
    .S(_0964_),
    .Z(_0966_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2456_ (.I(_0966_),
    .Z(_0175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2457_ (.A1(\wb_cross_clk.m_s_sync.s_data_ff[34] ),
    .A2(_0923_),
    .ZN(_0967_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2458_ (.A1(_0468_),
    .A2(_0925_),
    .B(_0967_),
    .ZN(_0176_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2459_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[35] ),
    .I1(_1567_),
    .S(_0964_),
    .Z(_0968_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2460_ (.I(_0968_),
    .Z(_0177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2461_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[36] ),
    .I1(_1560_),
    .S(_0964_),
    .Z(_0969_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2462_ (.I(_0969_),
    .Z(_0178_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2463_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[37] ),
    .I1(_1561_),
    .S(_0964_),
    .Z(_0970_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2464_ (.I(_0970_),
    .Z(_0179_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2465_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[38] ),
    .I1(_1574_),
    .S(_0964_),
    .Z(_0971_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2466_ (.I(_0971_),
    .Z(_0180_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2467_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[39] ),
    .I1(_1584_),
    .S(_0964_),
    .Z(_0972_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2468_ (.I(_0972_),
    .Z(_0181_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2469_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[40] ),
    .I1(_1575_),
    .S(_0964_),
    .Z(_0973_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2470_ (.I(_0973_),
    .Z(_0182_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2471_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[41] ),
    .I1(_1583_),
    .S(_0964_),
    .Z(_0974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2472_ (.I(_0974_),
    .Z(_0183_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2473_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[42] ),
    .I1(_1579_),
    .S(_0964_),
    .Z(_0975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2474_ (.I(_0975_),
    .Z(_0184_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2475_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[43] ),
    .I1(_1572_),
    .S(_0885_),
    .Z(_0976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2476_ (.I(_0976_),
    .Z(_0185_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2477_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[44] ),
    .I1(_1571_),
    .S(_0885_),
    .Z(_0977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2478_ (.I(_0977_),
    .Z(_0186_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2479_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[45] ),
    .I1(_0391_),
    .S(_0885_),
    .Z(_0978_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2480_ (.I(_0978_),
    .Z(_0187_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2481_ (.I0(\wb_cross_clk.m_s_sync.s_data_ff[46] ),
    .I1(_0525_),
    .S(_0885_),
    .Z(_0979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2482_ (.I(_0979_),
    .Z(_0188_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2483_ (.A1(\wb_cross_clk.s_m_sync.s_xfer_xor_flag ),
    .A2(_0676_),
    .Z(_0980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2484_ (.A1(_0553_),
    .A2(_0980_),
    .ZN(_0189_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2485_ (.A1(\wb_cross_clk.s_m_sync.s_xfer_xor_flag ),
    .A2(_0623_),
    .Z(_0981_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2486_ (.I(_0981_),
    .Z(_0190_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2487_ (.A1(_0623_),
    .A2(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[0] ),
    .Z(_0982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2488_ (.I(_0982_),
    .Z(_0191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2489_ (.A1(_0623_),
    .A2(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[1] ),
    .Z(_0983_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2490_ (.I(_0983_),
    .Z(_0192_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2491_ (.A1(_0634_),
    .A2(_0880_),
    .ZN(_0193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2492_ (.A1(\wb_cross_clk.msy_xor_err ),
    .A2(_0623_),
    .Z(_0984_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2493_ (.I(_0984_),
    .Z(_0194_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2494_ (.A1(_0922_),
    .A2(net209),
    .Z(_0985_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2495_ (.A1(_0634_),
    .A2(_0985_),
    .ZN(_0195_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2496_ (.A1(\wb_cross_clk.m_burst_cnt[0] ),
    .A2(_0878_),
    .Z(_0986_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2497_ (.A1(\wb_cross_clk.m_burst_cnt[0] ),
    .A2(_0878_),
    .B(_0885_),
    .ZN(_0987_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2498_ (.I(_0524_),
    .Z(_0988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2499_ (.A1(_1527_),
    .A2(net1),
    .ZN(_0989_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2500_ (.A1(_0933_),
    .A2(net210),
    .ZN(_0990_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2501_ (.A1(_0926_),
    .A2(_0989_),
    .B(_0990_),
    .ZN(_0991_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2502_ (.A1(_0986_),
    .A2(_0987_),
    .B(_0988_),
    .C(_0991_),
    .ZN(_0196_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2503_ (.A1(\wb_cross_clk.m_burst_cnt[1] ),
    .A2(\wb_cross_clk.m_burst_cnt[0] ),
    .A3(_0878_),
    .Z(_0992_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2504_ (.A1(\wb_cross_clk.m_burst_cnt[0] ),
    .A2(_0878_),
    .B(\wb_cross_clk.m_burst_cnt[1] ),
    .ZN(_0993_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2505_ (.A1(_0992_),
    .A2(_0993_),
    .B(_0579_),
    .C(_0925_),
    .ZN(_0197_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2506_ (.A1(\wb_cross_clk.m_burst_cnt[2] ),
    .A2(_0992_),
    .Z(_0994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2507_ (.A1(_0933_),
    .A2(_0926_),
    .ZN(_0995_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2508_ (.A1(_0923_),
    .A2(_0994_),
    .B1(_0995_),
    .B2(_0928_),
    .ZN(_0996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2509_ (.A1(_0623_),
    .A2(_0996_),
    .Z(_0997_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2510_ (.I(_0997_),
    .Z(_0198_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2511_ (.A1(\wb_cross_clk.m_burst_cnt[2] ),
    .A2(_0992_),
    .ZN(_0998_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2512_ (.A1(\wb_cross_clk.m_burst_cnt[3] ),
    .A2(_0998_),
    .ZN(_0999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2513_ (.A1(_0926_),
    .A2(_0990_),
    .B1(_0999_),
    .B2(_0885_),
    .ZN(_1000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2514_ (.A1(_0623_),
    .A2(_1000_),
    .Z(_1001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2515_ (.I(_1001_),
    .Z(_0199_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2516_ (.A1(\wb_cross_clk.s_burst_cnt[2] ),
    .A2(\wb_cross_clk.s_burst_cnt[1] ),
    .A3(\wb_cross_clk.s_burst_cnt[0] ),
    .Z(_1002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2517_ (.A1(\wb_compressor.wb_ack ),
    .A2(\wb_compressor.wb_err ),
    .B1(\wb_cross_clk.s_burst_cnt[3] ),
    .B2(_1002_),
    .ZN(_1003_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2518_ (.A1(_0933_),
    .A2(net240),
    .Z(_1004_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2519_ (.A1(\wb_cross_clk.m_s_sync.d_data[0] ),
    .A2(\wb_cross_clk.prev_xor_newreq ),
    .Z(_1005_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2520_ (.A1(_0676_),
    .A2(_1005_),
    .ZN(_1006_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2521_ (.A1(net240),
    .A2(_1006_),
    .ZN(_1007_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2522_ (.A1(\wb_cross_clk.m_s_sync.d_data[2] ),
    .A2(\wb_cross_clk.m_s_sync.d_data[1] ),
    .B(_1004_),
    .C(_1007_),
    .ZN(_1008_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2523_ (.A1(net240),
    .A2(_1006_),
    .Z(_1009_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2524_ (.A1(\wb_cross_clk.s_burst_cnt[0] ),
    .A2(net240),
    .ZN(_1010_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2525_ (.A1(\wb_cross_clk.s_burst_cnt[0] ),
    .A2(_1009_),
    .B(_1010_),
    .ZN(_1011_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2526_ (.A1(_1008_),
    .A2(_1011_),
    .B(_0549_),
    .ZN(_0200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2527_ (.A1(\wb_cross_clk.s_burst_cnt[1] ),
    .A2(_1006_),
    .ZN(_1012_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2528_ (.I0(_1012_),
    .I1(\wb_cross_clk.s_burst_cnt[1] ),
    .S(_1010_),
    .Z(_1013_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2529_ (.A1(_1008_),
    .A2(_1013_),
    .B(_0549_),
    .ZN(_0201_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2530_ (.A1(\wb_cross_clk.s_burst_cnt[1] ),
    .A2(\wb_cross_clk.s_burst_cnt[0] ),
    .B(\wb_cross_clk.s_burst_cnt[2] ),
    .ZN(_1014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2531_ (.A1(_1002_),
    .A2(_1014_),
    .B(net240),
    .ZN(_1015_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2532_ (.A1(\wb_cross_clk.m_s_sync.d_data[1] ),
    .A2(_1004_),
    .B(_1009_),
    .C(_1015_),
    .ZN(_1016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2533_ (.A1(\wb_cross_clk.s_burst_cnt[2] ),
    .A2(_1007_),
    .ZN(_1017_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2534_ (.A1(_0543_),
    .A2(_1016_),
    .A3(_1017_),
    .ZN(_0202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2535_ (.A1(\wb_compressor.wb_ack ),
    .A2(\wb_compressor.wb_err ),
    .B(_1002_),
    .ZN(_1018_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2536_ (.I(\wb_cross_clk.s_burst_cnt[3] ),
    .ZN(_1019_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2537_ (.A1(_1018_),
    .A2(_1007_),
    .B(_1019_),
    .C(_0660_),
    .ZN(_0203_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2538_ (.A1(_0528_),
    .A2(_1005_),
    .B(_0676_),
    .ZN(_1020_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2539_ (.A1(net240),
    .A2(_1020_),
    .ZN(_1021_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2540_ (.A1(_0553_),
    .A2(_1021_),
    .ZN(_0204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2541_ (.A1(_0553_),
    .A2(_0680_),
    .ZN(_0205_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2542_ (.A1(_0553_),
    .A2(_0678_),
    .ZN(_0206_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2543_ (.A1(\wb_cross_clk.msy_xor_ack ),
    .A2(_0623_),
    .Z(_1022_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2544_ (.I(_1022_),
    .Z(_0207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2545_ (.A1(_0768_),
    .A2(_0544_),
    .ZN(_0208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2546_ (.A1(\wb_compressor.state[4] ),
    .A2(\wb_compressor.state[1] ),
    .Z(_1023_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2547_ (.A1(\wb_compressor.state[6] ),
    .A2(\wb_compressor.state[3] ),
    .A3(_1023_),
    .ZN(_1024_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2548_ (.A1(\wb_compressor.state[5] ),
    .A2(\wb_compressor.state[2] ),
    .ZN(_1025_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2549_ (.A1(_1024_),
    .A2(_1025_),
    .ZN(_1026_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2550_ (.A1(_0542_),
    .A2(_0575_),
    .A3(_1026_),
    .ZN(_1027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2551_ (.A1(\wb_cross_clk.m_s_sync.d_data[5] ),
    .A2(_0458_),
    .ZN(_1028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2552_ (.A1(_1554_),
    .A2(_0933_),
    .B(_1028_),
    .ZN(_1029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2553_ (.A1(_1027_),
    .A2(_1029_),
    .ZN(_1030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2554_ (.A1(_0546_),
    .A2(_1027_),
    .B(_1030_),
    .ZN(_0209_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2555_ (.A1(\wb_cross_clk.m_s_sync.d_data[1] ),
    .A2(_1553_),
    .ZN(_1031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2556_ (.A1(_0415_),
    .A2(_0926_),
    .B(_1031_),
    .ZN(_1032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2557_ (.I(_0559_),
    .Z(_1033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2558_ (.A1(\wb_cross_clk.m_s_sync.d_data[2] ),
    .A2(_1033_),
    .ZN(_1034_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2559_ (.A1(_1033_),
    .A2(_0989_),
    .B(_1032_),
    .C(_1034_),
    .ZN(_1035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2560_ (.A1(net487),
    .A2(net220),
    .B(_1027_),
    .ZN(_1036_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2561_ (.A1(_0535_),
    .A2(_1027_),
    .B(net488),
    .ZN(_0210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2562_ (.I0(\wb_compressor.burst_end[2] ),
    .I1(net487),
    .S(_1027_),
    .Z(_1037_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2563_ (.I(_1037_),
    .Z(_0211_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2564_ (.A1(_0542_),
    .A2(_0533_),
    .A3(_0662_),
    .ZN(_1038_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _2565_ (.I(net213),
    .Z(_1039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2566_ (.I0(\wb_compressor.wb_i_dat[0] ),
    .I1(net67),
    .S(_1039_),
    .Z(_1040_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2567_ (.I(_1040_),
    .Z(_0212_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2568_ (.I0(\wb_compressor.wb_i_dat[1] ),
    .I1(net68),
    .S(_1039_),
    .Z(_1041_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2569_ (.I(_1041_),
    .Z(_0213_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2570_ (.I0(\wb_compressor.wb_i_dat[2] ),
    .I1(net69),
    .S(_1039_),
    .Z(_1042_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2571_ (.I(_1042_),
    .Z(_0214_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2572_ (.I0(\wb_compressor.wb_i_dat[3] ),
    .I1(net70),
    .S(_1039_),
    .Z(_1043_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2573_ (.I(_1043_),
    .Z(_0215_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2574_ (.I0(\wb_compressor.wb_i_dat[4] ),
    .I1(net71),
    .S(_1039_),
    .Z(_1044_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2575_ (.I(_1044_),
    .Z(_0216_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2576_ (.I0(\wb_compressor.wb_i_dat[5] ),
    .I1(net72),
    .S(_1039_),
    .Z(_1045_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2577_ (.I(_1045_),
    .Z(_0217_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2578_ (.I0(\wb_compressor.wb_i_dat[6] ),
    .I1(net73),
    .S(_1039_),
    .Z(_1046_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2579_ (.I(_1046_),
    .Z(_0218_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2580_ (.I0(\wb_compressor.wb_i_dat[7] ),
    .I1(net74),
    .S(_1039_),
    .Z(_1047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2581_ (.I(_1047_),
    .Z(_0219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2582_ (.I0(\wb_compressor.wb_i_dat[8] ),
    .I1(net75),
    .S(_1039_),
    .Z(_1048_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2583_ (.I(_1048_),
    .Z(_0220_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2584_ (.I0(\wb_compressor.wb_i_dat[9] ),
    .I1(net76),
    .S(_1039_),
    .Z(_1049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2585_ (.I(_1049_),
    .Z(_0221_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2586_ (.I0(\wb_compressor.wb_i_dat[10] ),
    .I1(net78),
    .S(net213),
    .Z(_1050_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2587_ (.I(_1050_),
    .Z(_0222_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2588_ (.I0(\wb_compressor.wb_i_dat[11] ),
    .I1(net79),
    .S(net212),
    .Z(_1051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2589_ (.I(_1051_),
    .Z(_0223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2590_ (.I0(\wb_compressor.wb_i_dat[12] ),
    .I1(net80),
    .S(net212),
    .Z(_1052_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2591_ (.I(_1052_),
    .Z(_0224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2592_ (.I0(\wb_compressor.wb_i_dat[13] ),
    .I1(net81),
    .S(net212),
    .Z(_1053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2593_ (.I(_1053_),
    .Z(_0225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2594_ (.I0(\wb_compressor.wb_i_dat[14] ),
    .I1(net82),
    .S(net214),
    .Z(_1054_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2595_ (.I(_1054_),
    .Z(_0226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2596_ (.I0(\wb_compressor.wb_i_dat[15] ),
    .I1(net83),
    .S(net214),
    .Z(_1055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2597_ (.I(_1055_),
    .Z(_0227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2598_ (.A1(\wb_compressor.wb_err ),
    .A2(_0662_),
    .B1(_0669_),
    .B2(net85),
    .ZN(_1056_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2599_ (.A1(\wb_compressor.state[1] ),
    .A2(\wb_compressor.state[6] ),
    .A3(_0543_),
    .A4(_1056_),
    .ZN(_1057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2600_ (.I(_1057_),
    .Z(_0228_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2601_ (.A1(\wb_compressor.wb_ack ),
    .A2(_0662_),
    .B1(_0669_),
    .B2(net84),
    .ZN(_1058_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2602_ (.A1(\wb_compressor.state[1] ),
    .A2(\wb_compressor.state[6] ),
    .A3(_0543_),
    .A4(_1058_),
    .ZN(_1059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2603_ (.I(_1059_),
    .Z(_0229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2604_ (.A1(_0641_),
    .A2(net91),
    .Z(_1060_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2605_ (.I(_1060_),
    .Z(_0230_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2606_ (.A1(_0641_),
    .A2(\sspi.sy_clk[0] ),
    .Z(_1061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2607_ (.I(_1061_),
    .Z(_0231_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2608_ (.A1(_0641_),
    .A2(\sspi.sy_clk[1] ),
    .Z(_1062_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2609_ (.I(_1062_),
    .Z(_0232_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2610_ (.A1(_0634_),
    .A2(_0581_),
    .ZN(_0233_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2611_ (.A1(\wb_compressor.state[1] ),
    .A2(\wb_compressor.state[6] ),
    .A3(_0665_),
    .B(_0666_),
    .ZN(_1063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2612_ (.A1(net250),
    .A2(_1063_),
    .ZN(_1064_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2613_ (.A1(net250),
    .A2(_0533_),
    .A3(_0540_),
    .B(_0545_),
    .ZN(_1065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2614_ (.A1(\wb_compressor.state[5] ),
    .A2(\wb_compressor.state[4] ),
    .B(_0666_),
    .C(_1065_),
    .ZN(_1066_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2615_ (.A1(_1064_),
    .A2(_1066_),
    .B(_0549_),
    .ZN(_0234_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2616_ (.A1(_0575_),
    .A2(_1024_),
    .ZN(_1067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2617_ (.A1(_1025_),
    .A2(_1067_),
    .B(net202),
    .ZN(_1068_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2618_ (.A1(\wb_compressor.state[5] ),
    .A2(\wb_compressor.state[2] ),
    .A3(_0551_),
    .A4(_1024_),
    .ZN(_1069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2619_ (.A1(_0543_),
    .A2(_1068_),
    .A3(_1069_),
    .ZN(_0235_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2620_ (.I(_1026_),
    .ZN(_1070_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2621_ (.A1(\wb_compressor.state[6] ),
    .A2(_0531_),
    .B1(_0575_),
    .B2(_1070_),
    .C(_1023_),
    .ZN(_1071_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2622_ (.I(net206),
    .Z(_1072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2623_ (.I(_1554_),
    .Z(_1073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2624_ (.I(_0458_),
    .Z(_1074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2625_ (.A1(\wb_cross_clk.m_s_sync.d_data[22] ),
    .A2(_1074_),
    .ZN(_1075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2626_ (.A1(_1073_),
    .A2(_0463_),
    .B(_1075_),
    .ZN(_1076_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2627_ (.A1(_0550_),
    .A2(_1025_),
    .ZN(_1077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2628_ (.A1(_0555_),
    .A2(_1077_),
    .ZN(_1078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2629_ (.I(_1078_),
    .Z(_1079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2630_ (.I(_1033_),
    .Z(_1080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2631_ (.A1(\wb_cross_clk.m_s_sync.d_data[6] ),
    .A2(_1080_),
    .B(_1077_),
    .ZN(_1081_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2632_ (.A1(_1080_),
    .A2(_1552_),
    .B(_1081_),
    .ZN(_1082_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2633_ (.A1(_0556_),
    .A2(_1076_),
    .B(_1079_),
    .C(_1082_),
    .ZN(_1083_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2634_ (.I(net206),
    .Z(_1084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2635_ (.A1(net176),
    .A2(_1084_),
    .ZN(_1085_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2636_ (.A1(_1072_),
    .A2(_1083_),
    .B(_1085_),
    .C(_0660_),
    .ZN(_0236_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2637_ (.I(_1077_),
    .Z(_1086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2638_ (.A1(net141),
    .A2(_1086_),
    .B1(_1079_),
    .B2(_0929_),
    .ZN(_1087_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2639_ (.A1(\wb_cross_clk.m_s_sync.d_data[23] ),
    .A2(_0458_),
    .ZN(_1088_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2640_ (.A1(_1554_),
    .A2(_0408_),
    .B(_1088_),
    .ZN(_1089_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2641_ (.A1(\wb_cross_clk.m_s_sync.d_data[7] ),
    .A2(_1077_),
    .B1(_1078_),
    .B2(\wb_cross_clk.m_s_sync.d_data[3] ),
    .ZN(_1090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2642_ (.I(_1090_),
    .ZN(_1091_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2643_ (.A1(_0555_),
    .A2(_1089_),
    .B1(_1091_),
    .B2(_1074_),
    .ZN(_1092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2644_ (.I(net207),
    .Z(_1093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2645_ (.A1(_1073_),
    .A2(_1087_),
    .B(_1092_),
    .C(_1093_),
    .ZN(_1094_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2646_ (.A1(net177),
    .A2(_1072_),
    .B(_1094_),
    .ZN(_1095_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2647_ (.A1(_0553_),
    .A2(_1095_),
    .ZN(_0237_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2648_ (.A1(net142),
    .A2(_1086_),
    .B1(_1079_),
    .B2(_0931_),
    .ZN(_1096_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2649_ (.I0(\wb_cross_clk.m_s_sync.d_data[24] ),
    .I1(net534),
    .S(_0559_),
    .Z(_1097_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2650_ (.A1(\wb_cross_clk.m_s_sync.d_data[8] ),
    .A2(_1077_),
    .B1(_1078_),
    .B2(\wb_cross_clk.m_s_sync.d_data[4] ),
    .ZN(_1098_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2651_ (.I(_1098_),
    .ZN(_1099_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2652_ (.A1(_0555_),
    .A2(_1097_),
    .B1(_1099_),
    .B2(_1074_),
    .ZN(_1100_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2653_ (.A1(_1073_),
    .A2(_1096_),
    .B(_1100_),
    .C(_1093_),
    .ZN(_1101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2654_ (.A1(net178),
    .A2(_1072_),
    .B(_1101_),
    .ZN(_1102_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2655_ (.A1(_0553_),
    .A2(_1102_),
    .ZN(_0238_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2656_ (.A1(_1073_),
    .A2(net528),
    .ZN(_1103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2657_ (.A1(\wb_cross_clk.m_s_sync.d_data[25] ),
    .A2(_1080_),
    .B(_0556_),
    .ZN(_1104_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2658_ (.A1(\wb_cross_clk.m_s_sync.d_data[9] ),
    .A2(_0428_),
    .ZN(_1105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2659_ (.A1(_1554_),
    .A2(_1539_),
    .B(_1105_),
    .ZN(_1106_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2660_ (.A1(_1029_),
    .A2(_1079_),
    .B1(_1106_),
    .B2(_1086_),
    .ZN(_1107_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2661_ (.A1(_1103_),
    .A2(_1104_),
    .B(_1107_),
    .C(_1093_),
    .ZN(_1108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2662_ (.A1(net179),
    .A2(_1072_),
    .B(_1108_),
    .ZN(_1109_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2663_ (.A1(_0553_),
    .A2(_1109_),
    .ZN(_0239_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2664_ (.A1(_1033_),
    .A2(_1593_),
    .ZN(_1110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2665_ (.A1(\wb_cross_clk.m_s_sync.d_data[26] ),
    .A2(_1080_),
    .B(_0555_),
    .C(_1110_),
    .ZN(_1111_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2666_ (.A1(\wb_cross_clk.m_s_sync.d_data[10] ),
    .A2(_0428_),
    .ZN(_1112_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2667_ (.A1(_1074_),
    .A2(net234),
    .B(_1112_),
    .ZN(_1113_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2668_ (.A1(net487),
    .A2(_1079_),
    .B1(_1113_),
    .B2(_1086_),
    .ZN(_1114_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2669_ (.A1(_1093_),
    .A2(_1111_),
    .A3(_1114_),
    .ZN(_1115_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2670_ (.A1(net180),
    .A2(_1084_),
    .B(_1115_),
    .ZN(_1116_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2671_ (.A1(_0774_),
    .A2(_1116_),
    .ZN(_0240_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2672_ (.A1(_1033_),
    .A2(_0406_),
    .ZN(_1117_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2673_ (.A1(\wb_cross_clk.m_s_sync.d_data[27] ),
    .A2(_1080_),
    .B(_0555_),
    .C(_1117_),
    .ZN(_1118_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2674_ (.A1(\wb_cross_clk.m_s_sync.d_data[11] ),
    .A2(_0428_),
    .ZN(_1119_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2675_ (.A1(_1554_),
    .A2(net235),
    .B(_1119_),
    .ZN(_1120_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2676_ (.A1(net220),
    .A2(_1079_),
    .B1(_1120_),
    .B2(_1086_),
    .ZN(_1121_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2677_ (.A1(_1093_),
    .A2(_1118_),
    .A3(_1121_),
    .ZN(_1122_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2678_ (.A1(net181),
    .A2(_1084_),
    .B(_1122_),
    .ZN(_1123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2679_ (.A1(_0774_),
    .A2(_1123_),
    .ZN(_0241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2680_ (.A1(\wb_cross_clk.m_s_sync.d_data[12] ),
    .A2(_1074_),
    .ZN(_1124_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2681_ (.A1(_1073_),
    .A2(net236),
    .B(_1124_),
    .ZN(_1125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2682_ (.I0(\wb_cross_clk.m_s_sync.d_data[28] ),
    .I1(net504),
    .S(_1033_),
    .Z(_1126_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2683_ (.A1(_1086_),
    .A2(_1125_),
    .B1(_1126_),
    .B2(_0556_),
    .ZN(_1127_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2684_ (.A1(net182),
    .A2(_1084_),
    .ZN(_1128_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2685_ (.A1(_1072_),
    .A2(net505),
    .B(_1128_),
    .C(_0660_),
    .ZN(_0242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2686_ (.A1(\wb_cross_clk.m_s_sync.d_data[13] ),
    .A2(_1074_),
    .ZN(_1129_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2687_ (.A1(_1073_),
    .A2(net237),
    .B(_1129_),
    .ZN(_1130_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2688_ (.I0(\wb_cross_clk.m_s_sync.d_data[29] ),
    .I1(net493),
    .S(_1033_),
    .Z(_1131_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2689_ (.A1(_1086_),
    .A2(_1130_),
    .B1(_1131_),
    .B2(_0556_),
    .ZN(_1132_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2690_ (.A1(net183),
    .A2(_1084_),
    .ZN(_1133_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2691_ (.A1(_1072_),
    .A2(net494),
    .B(_1133_),
    .C(_0660_),
    .ZN(_0243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2692_ (.A1(_1073_),
    .A2(net501),
    .ZN(_1134_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2693_ (.A1(\wb_cross_clk.m_s_sync.d_data[30] ),
    .A2(_1080_),
    .B(_0556_),
    .ZN(_1135_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2694_ (.I0(\wb_cross_clk.m_s_sync.d_data[14] ),
    .I1(net148),
    .S(_1033_),
    .Z(_1136_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2695_ (.A1(_0564_),
    .A2(_1078_),
    .B1(_1136_),
    .B2(_1086_),
    .ZN(_1137_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2696_ (.A1(_1134_),
    .A2(_1135_),
    .B(_1137_),
    .C(_1093_),
    .ZN(_1138_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2697_ (.A1(net184),
    .A2(_1084_),
    .B(net502),
    .ZN(_1139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2698_ (.A1(_0774_),
    .A2(_1139_),
    .ZN(_0244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2699_ (.A1(_1073_),
    .A2(net512),
    .ZN(_1140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2700_ (.A1(\wb_cross_clk.m_s_sync.d_data[31] ),
    .A2(_1080_),
    .B(_0556_),
    .ZN(_1141_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2701_ (.I0(\wb_cross_clk.m_s_sync.d_data[15] ),
    .I1(net149),
    .S(_1033_),
    .Z(_1142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2702_ (.A1(_0569_),
    .A2(_1078_),
    .B1(_1142_),
    .B2(_1086_),
    .ZN(_1143_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2703_ (.A1(_1140_),
    .A2(_1141_),
    .B(_1143_),
    .C(_1093_),
    .ZN(_1144_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2704_ (.A1(net185),
    .A2(_1084_),
    .B(net513),
    .ZN(_1145_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2705_ (.A1(_0774_),
    .A2(_1145_),
    .ZN(_0245_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2706_ (.A1(_1073_),
    .A2(net509),
    .ZN(_1146_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2707_ (.A1(\wb_cross_clk.m_s_sync.d_data[32] ),
    .A2(_1080_),
    .B(_0555_),
    .ZN(_1147_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2708_ (.I0(\wb_cross_clk.m_s_sync.d_data[16] ),
    .I1(net135),
    .S(_0559_),
    .Z(_1148_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2709_ (.A1(_0566_),
    .A2(_1078_),
    .B1(_1148_),
    .B2(_1086_),
    .ZN(_1149_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2710_ (.A1(_1146_),
    .A2(_1147_),
    .B(_1149_),
    .C(net208),
    .ZN(_1150_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2711_ (.A1(net187),
    .A2(_1084_),
    .B(net510),
    .ZN(_1151_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2712_ (.A1(_0774_),
    .A2(_1151_),
    .ZN(_0246_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2713_ (.A1(_1073_),
    .A2(net515),
    .ZN(_1152_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2714_ (.A1(\wb_cross_clk.m_s_sync.d_data[33] ),
    .A2(_1080_),
    .B(_0555_),
    .ZN(_1153_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2715_ (.I0(\wb_cross_clk.m_s_sync.d_data[17] ),
    .I1(net136),
    .S(_0559_),
    .Z(_1154_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2716_ (.A1(_0560_),
    .A2(_1078_),
    .B1(_1154_),
    .B2(_1077_),
    .ZN(_1155_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2717_ (.A1(_1152_),
    .A2(_1153_),
    .B(_1155_),
    .C(_1071_),
    .ZN(_1156_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2718_ (.A1(net188),
    .A2(_1084_),
    .B(net516),
    .ZN(_1157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2719_ (.A1(_0774_),
    .A2(_1157_),
    .ZN(_0247_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2720_ (.A1(\wb_compressor.state[5] ),
    .A2(\wb_compressor.state[6] ),
    .A3(\wb_compressor.state[2] ),
    .ZN(_1158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2721_ (.A1(_1554_),
    .A2(net137),
    .ZN(_1159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2722_ (.A1(\wb_cross_clk.m_s_sync.d_data[18] ),
    .A2(_1033_),
    .ZN(_1160_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2723_ (.A1(_1074_),
    .A2(net496),
    .ZN(_1161_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2724_ (.A1(\wb_cross_clk.m_s_sync.d_data[34] ),
    .A2(_1080_),
    .B(_0555_),
    .ZN(_1162_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2725_ (.A1(_1158_),
    .A2(_1159_),
    .A3(_1160_),
    .B1(_1161_),
    .B2(_1162_),
    .ZN(_1163_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2726_ (.A1(_0565_),
    .A2(_1079_),
    .B(net497),
    .ZN(_1164_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2727_ (.A1(net189),
    .A2(_1084_),
    .ZN(_1165_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2728_ (.A1(_1072_),
    .A2(net498),
    .B(_1165_),
    .C(_0660_),
    .ZN(_0248_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2729_ (.A1(_1554_),
    .A2(net138),
    .ZN(_1166_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2730_ (.A1(_0818_),
    .A2(_1074_),
    .B(_1158_),
    .C(_1166_),
    .ZN(_1167_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2731_ (.A1(_0556_),
    .A2(_0561_),
    .B1(_0572_),
    .B2(_1079_),
    .C(_1167_),
    .ZN(_1168_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2732_ (.A1(net190),
    .A2(_1093_),
    .ZN(_1169_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2733_ (.A1(_1072_),
    .A2(net217),
    .B(_1169_),
    .C(_0660_),
    .ZN(_0249_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2734_ (.A1(_1554_),
    .A2(net139),
    .ZN(_1170_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2735_ (.A1(_0820_),
    .A2(_1074_),
    .B(_1158_),
    .C(_1170_),
    .ZN(_1171_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2736_ (.A1(_0556_),
    .A2(_0570_),
    .B1(_0571_),
    .B2(_1079_),
    .C(_1171_),
    .ZN(_1172_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2737_ (.A1(net191),
    .A2(_1093_),
    .ZN(_1173_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2738_ (.A1(_1072_),
    .A2(net216),
    .B(_1173_),
    .C(_0660_),
    .ZN(_0250_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2739_ (.A1(_1554_),
    .A2(net140),
    .ZN(_1174_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2740_ (.A1(_0822_),
    .A2(_1074_),
    .B(_1158_),
    .C(_1174_),
    .ZN(_1175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2741_ (.A1(_0556_),
    .A2(_0562_),
    .B1(_0567_),
    .B2(_1079_),
    .C(_1175_),
    .ZN(_1176_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2742_ (.A1(net192),
    .A2(_1093_),
    .ZN(_1177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2743_ (.A1(_1072_),
    .A2(net215),
    .B(_1177_),
    .C(_0660_),
    .ZN(_0251_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2744_ (.A1(\sspi.state[5] ),
    .A2(_0624_),
    .ZN(_1178_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2745_ (.A1(\sspi.state[1] ),
    .A2(_1178_),
    .ZN(_1179_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2746_ (.A1(\sspi.state[0] ),
    .A2(_0618_),
    .ZN(_1180_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2747_ (.A1(\sspi.state[6] ),
    .A2(\sspi.state[2] ),
    .A3(\sspi.state[4] ),
    .ZN(_1181_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2748_ (.A1(_1180_),
    .A2(_1181_),
    .ZN(_1182_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2749_ (.A1(net254),
    .A2(_1182_),
    .ZN(_1183_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2750_ (.A1(_0597_),
    .A2(_1183_),
    .Z(_1184_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2751_ (.A1(_1527_),
    .A2(_0590_),
    .Z(_1185_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2752_ (.A1(\sspi.resp_err ),
    .A2(_1184_),
    .ZN(_1186_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2753_ (.A1(_1184_),
    .A2(_1185_),
    .B(_1186_),
    .C(_0917_),
    .ZN(_0252_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2754_ (.A1(\sspi.state[1] ),
    .A2(\sspi.state[3] ),
    .ZN(_1187_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2755_ (.A1(\sspi.state[6] ),
    .A2(_0639_),
    .A3(_1187_),
    .ZN(_1188_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2756_ (.I(_1188_),
    .ZN(_1189_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2757_ (.A1(\sspi.state[1] ),
    .A2(\sspi.state[6] ),
    .ZN(_1190_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2758_ (.A1(\sspi.state[3] ),
    .A2(\sspi.state[7] ),
    .B(_0617_),
    .ZN(_1191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2759_ (.A1(_1190_),
    .A2(_1191_),
    .B(\sspi.state[2] ),
    .ZN(_1192_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2760_ (.A1(_0639_),
    .A2(_1192_),
    .B(_1180_),
    .ZN(_1193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2761_ (.I(net243),
    .ZN(_1194_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2762_ (.A1(_0597_),
    .A2(_1189_),
    .B(_1194_),
    .ZN(_1195_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2763_ (.A1(_0602_),
    .A2(net204),
    .ZN(_1196_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2764_ (.A1(net243),
    .A2(_1188_),
    .ZN(_1197_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2765_ (.A1(\sspi.bit_cnt[0] ),
    .A2(_1197_),
    .B(_0641_),
    .ZN(_1198_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2766_ (.A1(_1196_),
    .A2(_1198_),
    .ZN(_0253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2767_ (.A1(\sspi.bit_cnt[1] ),
    .A2(net204),
    .ZN(_1199_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2768_ (.A1(\sspi.bit_cnt[1] ),
    .A2(\sspi.bit_cnt[0] ),
    .ZN(_1200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2769_ (.A1(_1200_),
    .A2(_0607_),
    .A3(_1197_),
    .ZN(_1201_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2770_ (.A1(_1199_),
    .A2(_1201_),
    .B(_0895_),
    .ZN(_0254_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2771_ (.I(\sspi.bit_cnt[2] ),
    .Z(_1202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2772_ (.A1(_1202_),
    .A2(net243),
    .B(_0603_),
    .ZN(_1203_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2773_ (.A1(_1189_),
    .A2(_1203_),
    .Z(_1204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2774_ (.A1(_1195_),
    .A2(_1204_),
    .B(_1202_),
    .ZN(_1205_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2775_ (.A1(_0603_),
    .A2(_1204_),
    .ZN(_1206_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2776_ (.I(_0579_),
    .Z(_1207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2777_ (.A1(_1205_),
    .A2(_1206_),
    .B(_1207_),
    .ZN(_0255_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2778_ (.I(\sspi.bit_cnt[3] ),
    .Z(_1208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2779_ (.A1(_0610_),
    .A2(net259),
    .Z(_1209_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2780_ (.A1(_1200_),
    .A2(net256),
    .ZN(_1210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2781_ (.A1(_1208_),
    .A2(net243),
    .B(_1210_),
    .ZN(_1211_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2782_ (.A1(_0609_),
    .A2(_0606_),
    .B1(_0637_),
    .B2(_0639_),
    .C(_1188_),
    .ZN(_1212_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2783_ (.A1(_1208_),
    .A2(net204),
    .B1(_1211_),
    .B2(_1212_),
    .ZN(_1213_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2784_ (.A1(_0634_),
    .A2(_1213_),
    .ZN(_0256_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2785_ (.A1(_0639_),
    .A2(_0636_),
    .B(_1210_),
    .ZN(_1214_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2786_ (.A1(\sspi.state[6] ),
    .A2(_1187_),
    .B(_1214_),
    .ZN(_1215_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2787_ (.I(_1215_),
    .ZN(_1216_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2788_ (.A1(_1195_),
    .A2(_1216_),
    .B(\sspi.bit_cnt[4] ),
    .ZN(_1217_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2789_ (.A1(_0600_),
    .A2(_0613_),
    .ZN(_1218_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2790_ (.A1(_0600_),
    .A2(_1210_),
    .B1(_1218_),
    .B2(net243),
    .ZN(_1219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2791_ (.A1(_0639_),
    .A2(_1219_),
    .ZN(_1220_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2792_ (.A1(_1217_),
    .A2(_1220_),
    .B(_1207_),
    .ZN(_0257_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2793_ (.A1(\sspi.state[0] ),
    .A2(\sspi.state[2] ),
    .A3(_0639_),
    .ZN(_1221_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2794_ (.A1(_1178_),
    .A2(_1190_),
    .A3(_1221_),
    .Z(_1222_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _2795_ (.A1(_0582_),
    .A2(_0597_),
    .A3(_1222_),
    .Z(_1223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2796_ (.I(_1223_),
    .Z(_1224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2797_ (.A1(\sspi.res_data[0] ),
    .A2(_1224_),
    .ZN(_1225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2798_ (.A1(_0516_),
    .A2(_0520_),
    .A3(_1223_),
    .Z(_1226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2799_ (.A1(_0988_),
    .A2(_1225_),
    .A3(_1226_),
    .ZN(_0258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2800_ (.I(_1223_),
    .Z(_1227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2801_ (.A1(_0510_),
    .A2(_0514_),
    .A3(_1227_),
    .Z(_1228_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2802_ (.I(_1223_),
    .Z(_1229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2803_ (.A1(\sspi.res_data[1] ),
    .A2(_1229_),
    .B(_0641_),
    .ZN(_1230_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2804_ (.A1(_1228_),
    .A2(_1230_),
    .ZN(_0259_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2805_ (.A1(_0504_),
    .A2(_0508_),
    .A3(_1227_),
    .Z(_1231_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2806_ (.A1(\sspi.res_data[2] ),
    .A2(_1229_),
    .B(_0641_),
    .ZN(_1232_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2807_ (.A1(_1231_),
    .A2(_1232_),
    .ZN(_0260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2808_ (.A1(_0498_),
    .A2(_0502_),
    .A3(_1227_),
    .Z(_1233_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2809_ (.A1(\sspi.res_data[3] ),
    .A2(_1224_),
    .B(_0641_),
    .ZN(_1234_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2810_ (.A1(_1233_),
    .A2(_1234_),
    .ZN(_0261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2811_ (.A1(_0492_),
    .A2(_0496_),
    .A3(_1227_),
    .Z(_1235_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2812_ (.A1(\sspi.res_data[4] ),
    .A2(_1224_),
    .B(_0763_),
    .ZN(_1236_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2813_ (.A1(_1235_),
    .A2(_1236_),
    .ZN(_0262_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2814_ (.A1(_0486_),
    .A2(_0490_),
    .A3(_1227_),
    .Z(_1237_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2815_ (.A1(\sspi.res_data[5] ),
    .A2(_1224_),
    .B(_0763_),
    .ZN(_1238_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2816_ (.A1(_1237_),
    .A2(_1238_),
    .ZN(_0263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2817_ (.A1(_0480_),
    .A2(_0484_),
    .A3(_1227_),
    .Z(_1239_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2818_ (.A1(\sspi.res_data[6] ),
    .A2(_1224_),
    .B(_0763_),
    .ZN(_1240_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2819_ (.A1(_1239_),
    .A2(_1240_),
    .ZN(_0264_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2820_ (.A1(_0460_),
    .A2(_0478_),
    .A3(_1223_),
    .Z(_1241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2821_ (.A1(\sspi.res_data[7] ),
    .A2(_1224_),
    .B(_0763_),
    .ZN(_1242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2822_ (.A1(_1241_),
    .A2(_1242_),
    .ZN(_0265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2823_ (.I(net125),
    .ZN(_1243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2824_ (.A1(\sspi.res_data[8] ),
    .A2(_1224_),
    .ZN(_1244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2825_ (.A1(_1243_),
    .A2(_1229_),
    .B(_1244_),
    .C(_0917_),
    .ZN(_0266_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2826_ (.I(net126),
    .ZN(_1245_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2827_ (.A1(\sspi.res_data[9] ),
    .A2(_1224_),
    .ZN(_1246_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2828_ (.A1(_1245_),
    .A2(_1229_),
    .B(_1246_),
    .C(_0917_),
    .ZN(_0267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2829_ (.I(net112),
    .ZN(_1247_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2830_ (.A1(\sspi.res_data[10] ),
    .A2(_1224_),
    .ZN(_1248_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2831_ (.A1(_1247_),
    .A2(_1229_),
    .B(_1248_),
    .C(_0917_),
    .ZN(_0268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2832_ (.I(net113),
    .ZN(_1249_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2833_ (.A1(\sspi.res_data[11] ),
    .A2(_1224_),
    .ZN(_1250_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2834_ (.A1(_1249_),
    .A2(_1229_),
    .B(_1250_),
    .C(_0917_),
    .ZN(_0269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2835_ (.I(net114),
    .ZN(_1251_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2836_ (.A1(\sspi.res_data[12] ),
    .A2(_1227_),
    .ZN(_1252_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2837_ (.I(_0579_),
    .Z(_1253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2838_ (.A1(_1251_),
    .A2(_1229_),
    .B(_1252_),
    .C(_1253_),
    .ZN(_0270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2839_ (.I(net115),
    .ZN(_1254_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2840_ (.A1(\sspi.res_data[13] ),
    .A2(_1227_),
    .ZN(_1255_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2841_ (.A1(_1254_),
    .A2(_1229_),
    .B(_1255_),
    .C(_1253_),
    .ZN(_0271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2842_ (.I(net116),
    .ZN(_1256_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2843_ (.A1(\sspi.res_data[14] ),
    .A2(_1227_),
    .ZN(_1257_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2844_ (.A1(_1256_),
    .A2(_1229_),
    .B(_1257_),
    .C(_1253_),
    .ZN(_0272_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2845_ (.I(net117),
    .ZN(_1258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2846_ (.A1(\sspi.res_data[15] ),
    .A2(_1227_),
    .ZN(_1259_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2847_ (.A1(_1258_),
    .A2(_1229_),
    .B(_1259_),
    .C(_1253_),
    .ZN(_0273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _2848_ (.I(net92),
    .ZN(_1260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2849_ (.A1(\sspi.state[6] ),
    .A2(_0582_),
    .A3(_1221_),
    .ZN(_1261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2850_ (.A1(_0611_),
    .A2(_1261_),
    .ZN(_1262_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2851_ (.A1(\sspi.req_data[0] ),
    .A2(_1262_),
    .B(_0763_),
    .ZN(_1263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2852_ (.A1(_1260_),
    .A2(_1262_),
    .B(_1263_),
    .ZN(_0274_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2853_ (.A1(_0635_),
    .A2(_1261_),
    .ZN(_1264_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2854_ (.A1(_0601_),
    .A2(\sspi.bit_cnt[0] ),
    .ZN(_1265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2855_ (.A1(_0605_),
    .A2(_1265_),
    .ZN(_1266_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2856_ (.A1(_0629_),
    .A2(net239),
    .A3(net253),
    .ZN(_1267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2857_ (.A1(net239),
    .A2(net253),
    .ZN(_1268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2858_ (.A1(\sspi.req_data[1] ),
    .A2(_1268_),
    .ZN(_1269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2859_ (.A1(_1267_),
    .A2(_1269_),
    .B(_1207_),
    .ZN(_0275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2860_ (.A1(\sspi.bit_cnt[1] ),
    .A2(_0602_),
    .ZN(_1270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2861_ (.A1(_0605_),
    .A2(_1270_),
    .ZN(_1271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2862_ (.A1(_0629_),
    .A2(_0611_),
    .A3(net239),
    .A4(_1271_),
    .ZN(_1272_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2863_ (.A1(net239),
    .A2(_1271_),
    .ZN(_1273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2864_ (.A1(\sspi.req_data[2] ),
    .A2(_1273_),
    .ZN(_1274_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2865_ (.A1(_1272_),
    .A2(_1274_),
    .B(_1207_),
    .ZN(_0276_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2866_ (.A1(_1200_),
    .A2(_0605_),
    .ZN(_1275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2867_ (.A1(_0629_),
    .A2(net239),
    .A3(_1275_),
    .ZN(_1276_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2868_ (.A1(net239),
    .A2(_1275_),
    .ZN(_1277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2869_ (.A1(\sspi.req_data[3] ),
    .A2(_1277_),
    .ZN(_1278_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2870_ (.A1(_1276_),
    .A2(_1278_),
    .B(_1207_),
    .ZN(_0277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2871_ (.A1(_1202_),
    .A2(_0619_),
    .A3(_0604_),
    .A4(_1264_),
    .ZN(_1279_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2872_ (.A1(_1202_),
    .A2(_0604_),
    .A3(net239),
    .ZN(_1280_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2873_ (.A1(\sspi.req_data[4] ),
    .A2(_1280_),
    .ZN(_1281_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2874_ (.A1(_1279_),
    .A2(_1281_),
    .B(_1207_),
    .ZN(_0278_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2875_ (.A1(\sspi.bit_cnt[1] ),
    .A2(_0602_),
    .ZN(_1282_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2876_ (.A1(_1209_),
    .A2(_0635_),
    .ZN(_1283_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2877_ (.A1(_1282_),
    .A2(_1283_),
    .ZN(_1284_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2878_ (.A1(_1261_),
    .A2(_1284_),
    .ZN(_1285_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2879_ (.A1(\sspi.req_data[5] ),
    .A2(_1285_),
    .B(_0763_),
    .ZN(_1286_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2880_ (.A1(_1260_),
    .A2(_1285_),
    .B(_1286_),
    .ZN(_0279_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2881_ (.A1(net92),
    .A2(_0611_),
    .ZN(_1287_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2882_ (.A1(_0601_),
    .A2(\sspi.bit_cnt[0] ),
    .ZN(_1288_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2883_ (.A1(_1288_),
    .A2(_1283_),
    .ZN(_1289_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2884_ (.A1(_1261_),
    .A2(_1289_),
    .ZN(_1290_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2885_ (.A1(\sspi.req_data[6] ),
    .A2(_1290_),
    .B(_0763_),
    .ZN(_1291_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2886_ (.A1(_1287_),
    .A2(_1290_),
    .B(_1291_),
    .ZN(_0280_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2887_ (.A1(_0606_),
    .A2(_0636_),
    .A3(_1261_),
    .ZN(_1292_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2888_ (.A1(\sspi.req_data[7] ),
    .A2(_1292_),
    .B(_0622_),
    .ZN(_1293_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2889_ (.A1(_1260_),
    .A2(_1292_),
    .B(_1293_),
    .ZN(_0281_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2890_ (.A1(\sspi.state[6] ),
    .A2(_0582_),
    .A3(_1221_),
    .Z(_1294_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2891_ (.I(_1294_),
    .Z(_1295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2892_ (.A1(_0609_),
    .A2(_1202_),
    .A3(_0607_),
    .ZN(_1296_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2893_ (.A1(_1295_),
    .A2(_1296_),
    .B(\sspi.req_data[8] ),
    .ZN(_1297_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2894_ (.A1(\sspi.bit_cnt[3] ),
    .A2(_0610_),
    .A3(net259),
    .ZN(_1298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2895_ (.A1(_0619_),
    .A2(_1261_),
    .A3(_1298_),
    .ZN(_1299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2896_ (.A1(_0988_),
    .A2(_1297_),
    .A3(_1299_),
    .ZN(_0282_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2897_ (.A1(_0619_),
    .A2(_0636_),
    .A3(_1295_),
    .A4(_1266_),
    .ZN(_1300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2898_ (.A1(_1208_),
    .A2(_1266_),
    .ZN(_1301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2899_ (.A1(_1261_),
    .A2(_1301_),
    .B(\sspi.req_data[9] ),
    .ZN(_1302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2900_ (.A1(_1300_),
    .A2(_1302_),
    .B(_1207_),
    .ZN(_0283_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2901_ (.A1(_0605_),
    .A2(_0608_),
    .A3(_1270_),
    .A4(_1287_),
    .ZN(_1303_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2902_ (.A1(_1208_),
    .A2(_1295_),
    .A3(_1271_),
    .ZN(_1304_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2903_ (.A1(_1295_),
    .A2(_1303_),
    .B1(_1304_),
    .B2(\sspi.req_data[10] ),
    .ZN(_1305_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2904_ (.A1(_0634_),
    .A2(_1305_),
    .ZN(_0284_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2905_ (.A1(_0619_),
    .A2(_0636_),
    .A3(_1275_),
    .Z(_1306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2906_ (.A1(_1208_),
    .A2(_1294_),
    .A3(_1275_),
    .ZN(_1307_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2907_ (.A1(_1295_),
    .A2(_1306_),
    .B1(_1307_),
    .B2(\sspi.req_data[11] ),
    .ZN(_1308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2908_ (.A1(_0634_),
    .A2(_1308_),
    .ZN(_0285_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2909_ (.A1(_0609_),
    .A2(_0610_),
    .A3(_1260_),
    .A4(_0607_),
    .ZN(_1309_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2910_ (.A1(_1208_),
    .A2(_1202_),
    .A3(net259),
    .A4(_1294_),
    .ZN(_1310_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2911_ (.A1(_1295_),
    .A2(_1309_),
    .B1(_1310_),
    .B2(\sspi.req_data[12] ),
    .ZN(_1311_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2912_ (.A1(_0634_),
    .A2(_1311_),
    .ZN(_0286_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2913_ (.A1(_0605_),
    .A2(_0636_),
    .A3(_1282_),
    .ZN(_1312_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2914_ (.A1(_1260_),
    .A2(_1312_),
    .ZN(_1313_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2915_ (.A1(_1295_),
    .A2(_1313_),
    .ZN(_1314_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2916_ (.A1(_1261_),
    .A2(_1312_),
    .B(\sspi.req_data[13] ),
    .ZN(_1315_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2917_ (.A1(_1314_),
    .A2(_1315_),
    .B(_1207_),
    .ZN(_0287_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2918_ (.A1(_0605_),
    .A2(_0636_),
    .A3(_1288_),
    .ZN(_1316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2919_ (.A1(_1287_),
    .A2(_1316_),
    .ZN(_1317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2920_ (.A1(_1295_),
    .A2(_1317_),
    .ZN(_1318_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2921_ (.A1(_1261_),
    .A2(_1316_),
    .B(\sspi.req_data[14] ),
    .ZN(_1319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2922_ (.A1(_1318_),
    .A2(_1319_),
    .B(_1207_),
    .ZN(_0288_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2923_ (.A1(_0629_),
    .A2(_0613_),
    .A3(_1295_),
    .ZN(_1320_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2924_ (.A1(_0613_),
    .A2(_1295_),
    .ZN(_1321_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2925_ (.A1(\sspi.req_data[15] ),
    .A2(_1321_),
    .ZN(_1322_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2926_ (.A1(_1320_),
    .A2(_1322_),
    .B(_1207_),
    .ZN(_0289_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2927_ (.A1(_0639_),
    .A2(_1180_),
    .ZN(_1323_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2928_ (.A1(\sspi.bit_cnt[4] ),
    .A2(_0611_),
    .A3(_1323_),
    .ZN(_1324_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2929_ (.A1(\sspi.req_addr[0] ),
    .A2(_1324_),
    .B(_0622_),
    .ZN(_1325_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2930_ (.A1(_1260_),
    .A2(net238),
    .B(_1325_),
    .ZN(_0290_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2931_ (.A1(_0639_),
    .A2(_1180_),
    .Z(_1326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2932_ (.A1(_0612_),
    .A2(net253),
    .A3(_1326_),
    .ZN(_1327_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2933_ (.A1(_0600_),
    .A2(_0611_),
    .Z(_1328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2934_ (.A1(_1327_),
    .A2(net252),
    .B(\sspi.req_addr[1] ),
    .ZN(_1329_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2935_ (.A1(_1323_),
    .A2(_1328_),
    .ZN(_1330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2936_ (.I(_1330_),
    .Z(_1331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2937_ (.A1(\sspi.bit_cnt[4] ),
    .A2(_0611_),
    .B(net92),
    .ZN(_1332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2938_ (.A1(_1208_),
    .A2(_0605_),
    .A3(_1265_),
    .A4(_1332_),
    .ZN(_1333_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2939_ (.A1(_1331_),
    .A2(_1333_),
    .ZN(_1334_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2940_ (.I(_0579_),
    .Z(_1335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2941_ (.A1(_1329_),
    .A2(_1334_),
    .B(_1335_),
    .ZN(_0291_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2942_ (.I(_1330_),
    .Z(_1336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2943_ (.A1(\sspi.bit_cnt[3] ),
    .A2(_0605_),
    .A3(_1270_),
    .ZN(_1337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2944_ (.A1(_1336_),
    .A2(_1337_),
    .ZN(_1338_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2945_ (.A1(\sspi.req_addr[2] ),
    .A2(_1338_),
    .ZN(_1339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2946_ (.A1(_0629_),
    .A2(_1331_),
    .A3(_1337_),
    .ZN(_1340_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2947_ (.A1(_1339_),
    .A2(_1340_),
    .B(_1335_),
    .ZN(_0292_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2948_ (.A1(\sspi.bit_cnt[3] ),
    .A2(_1200_),
    .A3(_0605_),
    .ZN(_1341_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2949_ (.A1(_1336_),
    .A2(net251),
    .B(\sspi.req_addr[3] ),
    .ZN(_1342_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2950_ (.A1(_1336_),
    .A2(_1332_),
    .A3(net251),
    .Z(_1343_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2951_ (.A1(_0988_),
    .A2(_1342_),
    .A3(_1343_),
    .ZN(_0293_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2952_ (.A1(\sspi.bit_cnt[3] ),
    .A2(_0610_),
    .A3(_0607_),
    .ZN(_1344_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2953_ (.A1(_1330_),
    .A2(_1344_),
    .ZN(_1345_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2954_ (.I0(_0619_),
    .I1(\sspi.req_addr[4] ),
    .S(_1345_),
    .Z(_1346_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2955_ (.A1(_0641_),
    .A2(_1346_),
    .Z(_1347_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2956_ (.I(_1347_),
    .Z(_0294_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2957_ (.A1(_1284_),
    .A2(_1332_),
    .ZN(_1348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2958_ (.A1(_1331_),
    .A2(_1348_),
    .ZN(_1349_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2959_ (.A1(\sspi.bit_cnt[4] ),
    .A2(_0611_),
    .Z(_1350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2960_ (.A1(_1326_),
    .A2(_1350_),
    .ZN(_1351_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2961_ (.A1(_1284_),
    .A2(_1351_),
    .B(\sspi.req_addr[5] ),
    .ZN(_1352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2962_ (.A1(_1349_),
    .A2(_1352_),
    .B(_1335_),
    .ZN(_0295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2963_ (.A1(_1289_),
    .A2(_1351_),
    .B(\sspi.req_addr[6] ),
    .ZN(_1353_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2964_ (.A1(net257),
    .A2(_0636_),
    .A3(_1270_),
    .ZN(_1354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2965_ (.A1(_0629_),
    .A2(_1354_),
    .A3(_1331_),
    .ZN(_1355_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2966_ (.A1(_1353_),
    .A2(_1355_),
    .B(_1335_),
    .ZN(_0296_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2967_ (.A1(_0606_),
    .A2(_0636_),
    .A3(_1332_),
    .ZN(_1356_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2968_ (.A1(_1210_),
    .A2(_0612_),
    .A3(_1336_),
    .ZN(_1357_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2969_ (.A1(_1331_),
    .A2(_1356_),
    .B1(_1357_),
    .B2(\sspi.req_addr[7] ),
    .ZN(_1358_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2970_ (.A1(_0580_),
    .A2(_1358_),
    .ZN(_0297_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2971_ (.A1(_1296_),
    .A2(_1336_),
    .B(\sspi.req_addr[8] ),
    .ZN(_1359_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2972_ (.A1(_0619_),
    .A2(_1298_),
    .A3(_1351_),
    .ZN(_1360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2973_ (.A1(_0988_),
    .A2(_1359_),
    .A3(_1360_),
    .ZN(_0298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2974_ (.A1(_0619_),
    .A2(_0636_),
    .A3(_1266_),
    .A4(_1336_),
    .ZN(_1361_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2975_ (.A1(_1301_),
    .A2(_1351_),
    .B(\sspi.req_addr[9] ),
    .ZN(_1362_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2976_ (.A1(_1361_),
    .A2(_1362_),
    .B(_1335_),
    .ZN(_0299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2977_ (.A1(_1208_),
    .A2(_1271_),
    .A3(_1336_),
    .ZN(_1363_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2978_ (.A1(_1303_),
    .A2(_1331_),
    .B1(_1363_),
    .B2(\sspi.req_addr[10] ),
    .ZN(_1364_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2979_ (.A1(_0580_),
    .A2(_1364_),
    .ZN(_0300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2980_ (.A1(_1208_),
    .A2(_1275_),
    .A3(_1336_),
    .ZN(_1365_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2981_ (.A1(_1306_),
    .A2(_1331_),
    .B1(_1365_),
    .B2(\sspi.req_addr[11] ),
    .ZN(_1366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2982_ (.A1(_0580_),
    .A2(_1366_),
    .ZN(_0301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2983_ (.A1(_1208_),
    .A2(_1202_),
    .A3(net259),
    .A4(_1336_),
    .ZN(_1367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2984_ (.A1(_1309_),
    .A2(_1331_),
    .B1(_1367_),
    .B2(\sspi.req_addr[12] ),
    .ZN(_1368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2985_ (.A1(_0580_),
    .A2(_1368_),
    .ZN(_0302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2986_ (.A1(_1313_),
    .A2(_1331_),
    .ZN(_1369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2987_ (.A1(_1312_),
    .A2(_1351_),
    .B(\sspi.req_addr[13] ),
    .ZN(_1370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2988_ (.A1(_1369_),
    .A2(_1370_),
    .B(_1335_),
    .ZN(_0303_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2989_ (.A1(_1317_),
    .A2(_1331_),
    .ZN(_1371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2990_ (.A1(_1316_),
    .A2(_1351_),
    .B(\sspi.req_addr[14] ),
    .ZN(_1372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2991_ (.A1(_1371_),
    .A2(_1372_),
    .B(_1335_),
    .ZN(_0304_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2992_ (.A1(_0629_),
    .A2(_0613_),
    .A3(_1336_),
    .ZN(_1373_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2993_ (.A1(_1218_),
    .A2(_1323_),
    .B(\sspi.req_addr[15] ),
    .ZN(_1374_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2994_ (.A1(_1373_),
    .A2(_1374_),
    .B(_1335_),
    .ZN(_0305_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2995_ (.A1(_0611_),
    .A2(_1323_),
    .ZN(_1375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2996_ (.I(_1332_),
    .ZN(_1376_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2997_ (.A1(\sspi.bit_cnt[4] ),
    .A2(_1375_),
    .ZN(_1377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2998_ (.A1(_1375_),
    .A2(_1376_),
    .B1(_1377_),
    .B2(\sspi.req_addr[16] ),
    .ZN(_1378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2999_ (.A1(_0580_),
    .A2(_1378_),
    .ZN(_0306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3000_ (.A1(_1327_),
    .A2(_1350_),
    .B(\sspi.req_addr[17] ),
    .ZN(_1379_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3001_ (.A1(_1323_),
    .A2(_1350_),
    .ZN(_1380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3002_ (.A1(_1333_),
    .A2(_1380_),
    .ZN(_1381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3003_ (.A1(_1379_),
    .A2(_1381_),
    .B(_1335_),
    .ZN(_0307_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3004_ (.I(\sspi.req_addr[18] ),
    .ZN(_1382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3005_ (.A1(_1337_),
    .A2(_1380_),
    .ZN(_1383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3006_ (.A1(_0629_),
    .A2(_1383_),
    .B(_0622_),
    .ZN(_1384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3007_ (.A1(_1382_),
    .A2(_1383_),
    .B(_1384_),
    .ZN(_0308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3008_ (.A1(net251),
    .A2(_1380_),
    .B(\sspi.req_addr[19] ),
    .ZN(_1385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3009_ (.A1(_1332_),
    .A2(net251),
    .A3(_1380_),
    .Z(_1386_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3010_ (.A1(_0988_),
    .A2(_1385_),
    .A3(_1386_),
    .ZN(_0309_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3011_ (.I(\sspi.req_addr[20] ),
    .ZN(_1387_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3012_ (.A1(_1344_),
    .A2(_1380_),
    .ZN(_1388_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3013_ (.A1(_0629_),
    .A2(_1388_),
    .B(_0622_),
    .ZN(_1389_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3014_ (.A1(_1387_),
    .A2(_1388_),
    .B(_1389_),
    .ZN(_0310_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3015_ (.A1(_1348_),
    .A2(_1380_),
    .ZN(_1390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3016_ (.A1(_1326_),
    .A2(net252),
    .ZN(_1391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3017_ (.A1(_1284_),
    .A2(_1391_),
    .B(\sspi.req_addr[21] ),
    .ZN(_1392_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3018_ (.A1(_1390_),
    .A2(_1392_),
    .B(_1335_),
    .ZN(_0311_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3019_ (.A1(_1354_),
    .A2(_1380_),
    .B(\sspi.req_addr[22] ),
    .ZN(_1393_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3020_ (.A1(_0619_),
    .A2(_1289_),
    .A3(_1391_),
    .ZN(_1394_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3021_ (.A1(_0988_),
    .A2(_1393_),
    .A3(_1394_),
    .ZN(_0312_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3022_ (.A1(net230),
    .A2(_1326_),
    .ZN(_1395_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3023_ (.A1(_1356_),
    .A2(_1380_),
    .B1(_1395_),
    .B2(\sspi.req_addr[23] ),
    .ZN(_1396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3024_ (.A1(_0580_),
    .A2(_1396_),
    .ZN(_0313_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3025_ (.I(\m_arbiter.wb0_we ),
    .ZN(_1397_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3026_ (.A1(_0524_),
    .A2(net254),
    .A3(_1182_),
    .ZN(_1398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3027_ (.I(_1398_),
    .Z(_1399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3028_ (.I(_1399_),
    .Z(_1400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3029_ (.A1(\sspi.state[1] ),
    .A2(_1399_),
    .ZN(_1401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3030_ (.I(_1401_),
    .Z(_1402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3031_ (.A1(_1397_),
    .A2(_1400_),
    .B(_1402_),
    .ZN(_0314_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3032_ (.I0(\sspi.req_data[0] ),
    .I1(\m_arbiter.wb0_o_dat[0] ),
    .S(_1402_),
    .Z(_1403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3033_ (.I(_1403_),
    .Z(_0315_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3034_ (.I0(\sspi.req_data[1] ),
    .I1(\m_arbiter.wb0_o_dat[1] ),
    .S(_1402_),
    .Z(_1404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3035_ (.I(_1404_),
    .Z(_0316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3036_ (.I0(\sspi.req_data[2] ),
    .I1(\m_arbiter.wb0_o_dat[2] ),
    .S(_1402_),
    .Z(_1405_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3037_ (.I(_1405_),
    .Z(_0317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3038_ (.I0(\sspi.req_data[3] ),
    .I1(\m_arbiter.wb0_o_dat[3] ),
    .S(_1402_),
    .Z(_1406_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3039_ (.I(_1406_),
    .Z(_0318_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3040_ (.I0(\sspi.req_data[4] ),
    .I1(\m_arbiter.wb0_o_dat[4] ),
    .S(_1402_),
    .Z(_1407_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3041_ (.I(_1407_),
    .Z(_0319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3042_ (.I0(\sspi.req_data[5] ),
    .I1(\m_arbiter.wb0_o_dat[5] ),
    .S(_1402_),
    .Z(_1408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3043_ (.I(_1408_),
    .Z(_0320_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3044_ (.I0(\sspi.req_data[6] ),
    .I1(\m_arbiter.wb0_o_dat[6] ),
    .S(_1402_),
    .Z(_1409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3045_ (.I(_1409_),
    .Z(_0321_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3046_ (.I0(\sspi.req_data[7] ),
    .I1(\m_arbiter.wb0_o_dat[7] ),
    .S(_1402_),
    .Z(_1410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3047_ (.I(_1410_),
    .Z(_0322_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3048_ (.I0(\sspi.req_data[8] ),
    .I1(\m_arbiter.wb0_o_dat[8] ),
    .S(_1402_),
    .Z(_1411_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3049_ (.I(_1411_),
    .Z(_0323_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3050_ (.I0(\sspi.req_data[9] ),
    .I1(\m_arbiter.wb0_o_dat[9] ),
    .S(_1401_),
    .Z(_1412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3051_ (.I(_1412_),
    .Z(_0324_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3052_ (.I0(\sspi.req_data[10] ),
    .I1(\m_arbiter.wb0_o_dat[10] ),
    .S(_1401_),
    .Z(_1413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3053_ (.I(_1413_),
    .Z(_0325_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3054_ (.I0(\sspi.req_data[11] ),
    .I1(\m_arbiter.wb0_o_dat[11] ),
    .S(_1401_),
    .Z(_1414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3055_ (.I(_1414_),
    .Z(_0326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3056_ (.I0(\sspi.req_data[12] ),
    .I1(\m_arbiter.wb0_o_dat[12] ),
    .S(_1401_),
    .Z(_1415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3057_ (.I(_1415_),
    .Z(_0327_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3058_ (.I0(\sspi.req_data[13] ),
    .I1(\m_arbiter.wb0_o_dat[13] ),
    .S(_1401_),
    .Z(_1416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3059_ (.I(_1416_),
    .Z(_0328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3060_ (.I0(\sspi.req_data[14] ),
    .I1(\m_arbiter.wb0_o_dat[14] ),
    .S(_1401_),
    .Z(_1417_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3061_ (.I(_1417_),
    .Z(_0329_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3062_ (.I0(\sspi.req_data[15] ),
    .I1(\m_arbiter.wb0_o_dat[15] ),
    .S(_1401_),
    .Z(_1418_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3063_ (.I(_1418_),
    .Z(_0330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3064_ (.I(net244),
    .Z(_1419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3065_ (.A1(\clk_div.cnt[0] ),
    .A2(_1419_),
    .ZN(_0331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3066_ (.A1(\clk_div.cnt[0] ),
    .A2(\clk_div.cnt[1] ),
    .ZN(_1420_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3067_ (.A1(_1419_),
    .A2(_1420_),
    .ZN(_0332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3068_ (.A1(\clk_div.cnt[0] ),
    .A2(\clk_div.cnt[1] ),
    .A3(\clk_div.cnt[2] ),
    .Z(_1421_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3069_ (.A1(\clk_div.cnt[0] ),
    .A2(\clk_div.cnt[1] ),
    .B(\clk_div.cnt[2] ),
    .ZN(_1422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3070_ (.A1(_1419_),
    .A2(_1421_),
    .A3(_1422_),
    .ZN(_0333_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _3071_ (.A1(\clk_div.cnt[0] ),
    .A2(\clk_div.cnt[1] ),
    .A3(\clk_div.cnt[2] ),
    .A4(\clk_div.cnt[3] ),
    .Z(_1423_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3072_ (.A1(\clk_div.cnt[3] ),
    .A2(_1421_),
    .ZN(_1424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3073_ (.A1(_1419_),
    .A2(_1423_),
    .A3(_1424_),
    .ZN(_0334_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3074_ (.A1(\clk_div.cnt[4] ),
    .A2(_1423_),
    .Z(_1425_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3075_ (.A1(_0756_),
    .A2(_1425_),
    .Z(_1426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3076_ (.I(_1426_),
    .Z(_0335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3077_ (.A1(\clk_div.cnt[4] ),
    .A2(_1423_),
    .ZN(_1427_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3078_ (.A1(\clk_div.cnt[5] ),
    .A2(_1427_),
    .Z(_1428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3079_ (.A1(_1419_),
    .A2(_1428_),
    .ZN(_0336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3080_ (.A1(\clk_div.cnt[4] ),
    .A2(\clk_div.cnt[5] ),
    .A3(_1423_),
    .ZN(_1429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3081_ (.A1(\clk_div.cnt[6] ),
    .A2(_1429_),
    .Z(_1430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3082_ (.A1(_1419_),
    .A2(_1430_),
    .ZN(_0337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3083_ (.I(\clk_div.cnt[7] ),
    .ZN(_1431_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3084_ (.A1(\clk_div.cnt[4] ),
    .A2(\clk_div.cnt[5] ),
    .A3(\clk_div.cnt[6] ),
    .A4(_1423_),
    .ZN(_1432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3085_ (.A1(_1431_),
    .A2(_1432_),
    .ZN(_1433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3086_ (.A1(_1431_),
    .A2(_1432_),
    .Z(_1434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3087_ (.A1(_1419_),
    .A2(_1433_),
    .A3(_1434_),
    .ZN(_0338_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3088_ (.I(\clk_div.cnt[8] ),
    .ZN(_1435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3089_ (.A1(_1431_),
    .A2(_1435_),
    .A3(_1432_),
    .ZN(_1436_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3090_ (.A1(\clk_div.cnt[8] ),
    .A2(_1433_),
    .ZN(_1437_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3091_ (.A1(_1419_),
    .A2(_1436_),
    .A3(_1437_),
    .ZN(_0339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3092_ (.A1(\clk_div.cnt[9] ),
    .A2(_1436_),
    .Z(_1438_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3093_ (.A1(\clk_div.cnt[9] ),
    .A2(_1436_),
    .ZN(_1439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3094_ (.A1(net244),
    .A2(_1438_),
    .A3(_1439_),
    .ZN(_0340_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3095_ (.A1(\clk_div.cnt[10] ),
    .A2(_1438_),
    .Z(_1440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3096_ (.A1(\clk_div.cnt[10] ),
    .A2(_1438_),
    .B(_0756_),
    .ZN(_1441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3097_ (.A1(_1440_),
    .A2(_1441_),
    .ZN(_0341_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3098_ (.A1(\clk_div.cnt[11] ),
    .A2(_1440_),
    .Z(_1442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3099_ (.A1(\clk_div.cnt[11] ),
    .A2(_1440_),
    .B(_0756_),
    .ZN(_1443_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3100_ (.A1(_1442_),
    .A2(_1443_),
    .ZN(_0342_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3101_ (.A1(\clk_div.cnt[12] ),
    .A2(_1442_),
    .Z(_1444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3102_ (.A1(\clk_div.cnt[12] ),
    .A2(_1442_),
    .B(_0756_),
    .ZN(_1445_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3103_ (.A1(_1444_),
    .A2(_1445_),
    .ZN(_0343_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3104_ (.A1(\clk_div.cnt[13] ),
    .A2(_1444_),
    .Z(_1446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3105_ (.A1(\clk_div.cnt[13] ),
    .A2(_1444_),
    .B(_0756_),
    .ZN(_1447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3106_ (.A1(_1446_),
    .A2(_1447_),
    .ZN(_0344_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3107_ (.A1(\clk_div.cnt[14] ),
    .A2(_1446_),
    .ZN(_1448_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3108_ (.A1(_1419_),
    .A2(_1448_),
    .ZN(_0345_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3109_ (.A1(\clk_div.cnt[14] ),
    .A2(_1446_),
    .B(\clk_div.cnt[15] ),
    .ZN(_1449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3110_ (.A1(_1419_),
    .A2(_1449_),
    .ZN(_0346_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3111_ (.A1(\m_arbiter.i_wb0_cyc ),
    .A2(_1183_),
    .B(_0763_),
    .ZN(_1450_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3112_ (.A1(_1184_),
    .A2(_1450_),
    .ZN(_0347_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3113_ (.A1(\sspi.state[5] ),
    .A2(\sspi.state[7] ),
    .ZN(_1451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3114_ (.A1(_1187_),
    .A2(_1451_),
    .ZN(_1452_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3115_ (.A1(net258),
    .A2(_1452_),
    .ZN(_1453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3116_ (.A1(_0621_),
    .A2(_1453_),
    .B(_0618_),
    .ZN(_1454_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3117_ (.A1(_0597_),
    .A2(_1179_),
    .B(_1454_),
    .ZN(_1455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3118_ (.A1(\sspi.res_data[3] ),
    .A2(_1200_),
    .B1(_1265_),
    .B2(\sspi.res_data[1] ),
    .ZN(_1456_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3119_ (.A1(\sspi.res_data[0] ),
    .A2(_0607_),
    .B1(_1270_),
    .B2(\sspi.res_data[2] ),
    .ZN(_1457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3120_ (.A1(_1202_),
    .A2(_1456_),
    .A3(_1457_),
    .ZN(_1458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3121_ (.A1(\sspi.res_data[4] ),
    .A2(net259),
    .B1(_1282_),
    .B2(\sspi.res_data[5] ),
    .ZN(_1459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3122_ (.A1(\sspi.res_data[7] ),
    .A2(_0603_),
    .B1(_1288_),
    .B2(\sspi.res_data[6] ),
    .ZN(_1460_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3123_ (.A1(_1459_),
    .A2(_1460_),
    .B(_0610_),
    .ZN(_1461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3124_ (.A1(\sspi.res_data[11] ),
    .A2(_0603_),
    .B1(_1288_),
    .B2(\sspi.res_data[10] ),
    .ZN(_1462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3125_ (.A1(\sspi.res_data[8] ),
    .A2(net259),
    .B1(_1282_),
    .B2(\sspi.res_data[9] ),
    .ZN(_1463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3126_ (.A1(_1462_),
    .A2(_1463_),
    .B(_1202_),
    .ZN(_1464_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3127_ (.A1(\sspi.res_data[14] ),
    .A2(_1270_),
    .B(_1202_),
    .ZN(_1465_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _3128_ (.A1(\sspi.res_data[15] ),
    .A2(_1200_),
    .B1(_0607_),
    .B2(\sspi.res_data[12] ),
    .C1(_1265_),
    .C2(\sspi.res_data[13] ),
    .ZN(_1466_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3129_ (.A1(_1465_),
    .A2(_1466_),
    .B(\sspi.bit_cnt[3] ),
    .ZN(_1467_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3130_ (.A1(\sspi.bit_cnt[3] ),
    .A2(net242),
    .A3(_1461_),
    .B1(_1464_),
    .B2(_1467_),
    .ZN(_1468_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3131_ (.A1(\sspi.state[3] ),
    .A2(net492),
    .B(_0617_),
    .ZN(_1469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3132_ (.A1(\sspi.resp_err ),
    .A2(_0617_),
    .B(_1469_),
    .ZN(_1470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3133_ (.A1(\sspi.state[1] ),
    .A2(_1470_),
    .B(_0621_),
    .ZN(_1471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3134_ (.A1(net195),
    .A2(_1455_),
    .B1(_1471_),
    .B2(_1454_),
    .ZN(_1472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3135_ (.A1(_0761_),
    .A2(_1472_),
    .ZN(_0348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3136_ (.I0(\m_arbiter.wb0_adr[0] ),
    .I1(\sspi.req_addr[0] ),
    .S(_1400_),
    .Z(_1473_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3137_ (.I(_1473_),
    .Z(_0349_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3138_ (.I0(\m_arbiter.wb0_adr[1] ),
    .I1(\sspi.req_addr[1] ),
    .S(_1400_),
    .Z(_1474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3139_ (.I(_1474_),
    .Z(_0350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3140_ (.I0(\m_arbiter.wb0_adr[2] ),
    .I1(\sspi.req_addr[2] ),
    .S(_1400_),
    .Z(_1475_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3141_ (.I(_1475_),
    .Z(_0351_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3142_ (.I0(\m_arbiter.wb0_adr[3] ),
    .I1(\sspi.req_addr[3] ),
    .S(_1400_),
    .Z(_1476_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3143_ (.I(_1476_),
    .Z(_0352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3144_ (.I0(\m_arbiter.wb0_adr[4] ),
    .I1(\sspi.req_addr[4] ),
    .S(_1400_),
    .Z(_1477_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3145_ (.I(_1477_),
    .Z(_0353_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3146_ (.I(_1399_),
    .Z(_1478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3147_ (.I0(\m_arbiter.wb0_adr[5] ),
    .I1(\sspi.req_addr[5] ),
    .S(_1478_),
    .Z(_1479_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3148_ (.I(_1479_),
    .Z(_0354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3149_ (.I0(\m_arbiter.wb0_adr[6] ),
    .I1(\sspi.req_addr[6] ),
    .S(_1478_),
    .Z(_1480_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3150_ (.I(_1480_),
    .Z(_0355_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3151_ (.I0(\m_arbiter.wb0_adr[7] ),
    .I1(\sspi.req_addr[7] ),
    .S(_1478_),
    .Z(_1481_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3152_ (.I(_1481_),
    .Z(_0356_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3153_ (.A1(\sspi.req_addr[8] ),
    .A2(_1400_),
    .ZN(_1482_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3154_ (.A1(_1555_),
    .A2(_1400_),
    .B(_1482_),
    .ZN(_0357_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3155_ (.I0(\m_arbiter.wb0_adr[9] ),
    .I1(\sspi.req_addr[9] ),
    .S(_1478_),
    .Z(_1483_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3156_ (.I(_1483_),
    .Z(_0358_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3157_ (.I0(\m_arbiter.wb0_adr[10] ),
    .I1(\sspi.req_addr[10] ),
    .S(_1478_),
    .Z(_1484_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3158_ (.I(_1484_),
    .Z(_0359_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3159_ (.I0(\m_arbiter.wb0_adr[11] ),
    .I1(\sspi.req_addr[11] ),
    .S(_1478_),
    .Z(_1485_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3160_ (.I(_1485_),
    .Z(_0360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3161_ (.I0(\m_arbiter.wb0_adr[12] ),
    .I1(\sspi.req_addr[12] ),
    .S(_1478_),
    .Z(_1486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3162_ (.I(_1486_),
    .Z(_0361_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3163_ (.I0(\m_arbiter.wb0_adr[13] ),
    .I1(\sspi.req_addr[13] ),
    .S(_1478_),
    .Z(_1487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3164_ (.I(_1487_),
    .Z(_0362_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3165_ (.I0(\m_arbiter.wb0_adr[14] ),
    .I1(\sspi.req_addr[14] ),
    .S(_1478_),
    .Z(_1488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3166_ (.I(_1488_),
    .Z(_0363_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3167_ (.I0(\m_arbiter.wb0_adr[15] ),
    .I1(\sspi.req_addr[15] ),
    .S(_1478_),
    .Z(_1489_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3168_ (.I(_1489_),
    .Z(_0364_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3169_ (.I0(\m_arbiter.wb0_adr[16] ),
    .I1(\sspi.req_addr[16] ),
    .S(_1399_),
    .Z(_1490_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3170_ (.I(_1490_),
    .Z(_0365_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3171_ (.I0(\m_arbiter.wb0_adr[17] ),
    .I1(\sspi.req_addr[17] ),
    .S(_1399_),
    .Z(_1491_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3172_ (.I(_1491_),
    .Z(_0366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3173_ (.I0(\m_arbiter.wb0_adr[18] ),
    .I1(\sspi.req_addr[18] ),
    .S(_1399_),
    .Z(_1492_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3174_ (.I(_1492_),
    .Z(_0367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3175_ (.I0(\m_arbiter.wb0_adr[19] ),
    .I1(\sspi.req_addr[19] ),
    .S(_1399_),
    .Z(_1493_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3176_ (.I(_1493_),
    .Z(_0368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3177_ (.I0(\m_arbiter.wb0_adr[20] ),
    .I1(\sspi.req_addr[20] ),
    .S(_1399_),
    .Z(_1494_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3178_ (.I(_1494_),
    .Z(_0369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3179_ (.I0(\m_arbiter.wb0_adr[21] ),
    .I1(\sspi.req_addr[21] ),
    .S(_1399_),
    .Z(_1495_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3180_ (.I(_1495_),
    .Z(_0370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3181_ (.I0(\m_arbiter.wb0_adr[22] ),
    .I1(\sspi.req_addr[22] ),
    .S(_1399_),
    .Z(_1496_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3182_ (.I(_1496_),
    .Z(_0371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3183_ (.A1(\sspi.req_addr[23] ),
    .A2(_1400_),
    .ZN(_1497_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3184_ (.A1(_1577_),
    .A2(_1400_),
    .B(_1497_),
    .ZN(_0372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3185_ (.A1(net241),
    .A2(net232),
    .A3(_0466_),
    .A4(_0658_),
    .ZN(_1498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3186_ (.I(_1498_),
    .Z(_1499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3187_ (.A1(net151),
    .A2(_1499_),
    .ZN(_1500_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3188_ (.A1(_1552_),
    .A2(_1499_),
    .B(_1500_),
    .C(_0761_),
    .ZN(_0373_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3189_ (.A1(net162),
    .A2(_1499_),
    .ZN(_1501_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3190_ (.A1(_1548_),
    .A2(_1499_),
    .B(_1501_),
    .C(_0761_),
    .ZN(_0374_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3191_ (.A1(net169),
    .A2(_1498_),
    .ZN(_1502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3192_ (.A1(_1544_),
    .A2(_1499_),
    .B(_1502_),
    .C(_0761_),
    .ZN(_0375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3193_ (.A1(net170),
    .A2(_1498_),
    .ZN(_1503_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3194_ (.A1(_1539_),
    .A2(_1499_),
    .B(_1503_),
    .C(_0761_),
    .ZN(_0376_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3195_ (.A1(net171),
    .A2(_1498_),
    .ZN(_1504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3196_ (.A1(net234),
    .A2(_1499_),
    .B(_1504_),
    .C(_0761_),
    .ZN(_0377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3197_ (.A1(net172),
    .A2(_1498_),
    .ZN(_1505_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3198_ (.A1(net235),
    .A2(_1499_),
    .B(_1505_),
    .C(_0761_),
    .ZN(_0378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3199_ (.A1(net173),
    .A2(_1498_),
    .ZN(_1506_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3200_ (.A1(net236),
    .A2(_1499_),
    .B(_1506_),
    .C(_0761_),
    .ZN(_0379_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3201_ (.A1(net174),
    .A2(_1498_),
    .ZN(_1507_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3202_ (.A1(net237),
    .A2(_1499_),
    .B(_1507_),
    .C(_0623_),
    .ZN(_0380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _3203_ (.A1(net241),
    .A2(_0464_),
    .A3(net233),
    .A4(_0658_),
    .Z(_1508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3204_ (.I(_1508_),
    .Z(_1509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3205_ (.A1(net175),
    .A2(_1509_),
    .ZN(_1510_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3206_ (.A1(_1552_),
    .A2(_1509_),
    .B(_1510_),
    .C(_1253_),
    .ZN(_0381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3207_ (.A1(net186),
    .A2(_1509_),
    .ZN(_1511_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3208_ (.A1(_1548_),
    .A2(_1509_),
    .B(_1511_),
    .C(_1253_),
    .ZN(_0382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3209_ (.A1(net194),
    .A2(_1508_),
    .ZN(_1512_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3210_ (.A1(_1544_),
    .A2(_1509_),
    .B(_1512_),
    .C(_1253_),
    .ZN(_0383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3211_ (.A1(net197),
    .A2(_1508_),
    .ZN(_1513_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3212_ (.A1(_1539_),
    .A2(_1509_),
    .B(_1513_),
    .C(_1253_),
    .ZN(_0384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3213_ (.A1(net198),
    .A2(_1508_),
    .ZN(_1514_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3214_ (.A1(net234),
    .A2(_1509_),
    .B(_1514_),
    .C(_1253_),
    .ZN(_0385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3215_ (.A1(net199),
    .A2(_1508_),
    .ZN(_1515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3216_ (.A1(net235),
    .A2(_1509_),
    .B(_1515_),
    .C(_1253_),
    .ZN(_0386_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3217_ (.A1(net200),
    .A2(_1508_),
    .ZN(_1516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3218_ (.A1(net236),
    .A2(_1509_),
    .B(_1516_),
    .C(_0988_),
    .ZN(_0387_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3219_ (.A1(net201),
    .A2(_1508_),
    .ZN(_1517_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3220_ (.A1(net237),
    .A2(_1509_),
    .B(_1517_),
    .C(_0988_),
    .ZN(_0388_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3221_ (.I(net64),
    .Z(_1518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _3222_ (.I(net65),
    .ZN(_1519_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3223_ (.I(net98),
    .Z(_1520_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3224_ (.A1(_1518_),
    .A2(_1519_),
    .B(_1520_),
    .ZN(_0015_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3225_ (.A1(_1518_),
    .A2(_1519_),
    .B(_1520_),
    .ZN(_0016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3226_ (.A1(_1518_),
    .A2(_1519_),
    .B(_1520_),
    .ZN(_0017_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3227_ (.A1(_1518_),
    .A2(_1519_),
    .B(_1520_),
    .ZN(_0018_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3228_ (.A1(_1518_),
    .A2(_1519_),
    .B(_1520_),
    .ZN(_0019_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3229_ (.A1(_1518_),
    .A2(_1519_),
    .B(_1520_),
    .ZN(_0020_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3230_ (.A1(_1518_),
    .A2(_1519_),
    .B(_1520_),
    .ZN(_0021_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3231_ (.A1(_1518_),
    .A2(_1519_),
    .B(_1520_),
    .ZN(_0022_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3232_ (.A1(_1527_),
    .A2(net27),
    .ZN(_1521_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3233_ (.A1(\m_arbiter.i_wb0_cyc ),
    .A2(_0523_),
    .B(_1521_),
    .C(_0988_),
    .ZN(_0389_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3234_ (.D(_0023_),
    .CLK(clknet_4_2_0_net196),
    .Q(\wb_compressor.burst_cnt[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3235_ (.D(_0024_),
    .CLK(clknet_4_0_0_net196),
    .Q(\wb_compressor.burst_cnt[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3236_ (.D(_0025_),
    .CLK(clknet_4_0_0_net196),
    .Q(\wb_compressor.burst_cnt[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3237_ (.D(net90),
    .CLK(clknet_leaf_3_user_clock2),
    .Q(\embed_s_ff[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3238_ (.D(net529),
    .CLK(clknet_leaf_13_user_clock2),
    .Q(net106),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3239_ (.D(net89),
    .CLK(clknet_leaf_3_user_clock2),
    .Q(\disable_s_ff[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3240_ (.D(net530),
    .CLK(clknet_leaf_13_user_clock2),
    .Q(net105),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3241_ (.D(net88),
    .CLK(clknet_leaf_0_user_clock2),
    .Q(\split_s_ff[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3242_ (.D(net532),
    .CLK(clknet_leaf_0_user_clock2),
    .Q(\clk_div.clock_sel ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3243_ (.D(net87),
    .CLK(clknet_leaf_13_user_clock2),
    .Q(\irq_s_ff[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3244_ (.D(net535),
    .CLK(clknet_leaf_13_user_clock2),
    .Q(net107),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3245_ (.D(_0026_),
    .CLK(clknet_4_14_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3246_ (.D(_0027_),
    .CLK(clknet_4_12_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3247_ (.D(_0028_),
    .CLK(clknet_4_14_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3248_ (.D(_0029_),
    .CLK(clknet_4_15_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3249_ (.D(_0030_),
    .CLK(clknet_4_15_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3250_ (.D(_0031_),
    .CLK(clknet_4_11_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3251_ (.D(_0032_),
    .CLK(clknet_4_15_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3252_ (.D(_0033_),
    .CLK(clknet_4_15_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3253_ (.D(_0034_),
    .CLK(clknet_4_13_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3254_ (.D(_0035_),
    .CLK(clknet_4_13_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3255_ (.D(_0036_),
    .CLK(clknet_4_15_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3256_ (.D(_0037_),
    .CLK(clknet_4_13_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3257_ (.D(_0038_),
    .CLK(clknet_4_5_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3258_ (.D(_0039_),
    .CLK(clknet_4_7_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3259_ (.D(_0040_),
    .CLK(clknet_4_5_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3260_ (.D(_0041_),
    .CLK(clknet_4_4_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3261_ (.D(_0042_),
    .CLK(clknet_4_7_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[16] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3262_ (.D(_0043_),
    .CLK(clknet_4_13_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[17] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3263_ (.D(_0044_),
    .CLK(clknet_leaf_31_user_clock2),
    .Q(iram_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3264_ (.D(_0045_),
    .CLK(clknet_leaf_30_user_clock2),
    .Q(\iram_latched[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3265_ (.D(_0046_),
    .CLK(clknet_leaf_30_user_clock2),
    .Q(\iram_latched[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3266_ (.D(_0047_),
    .CLK(clknet_leaf_30_user_clock2),
    .Q(\iram_latched[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3267_ (.D(_0048_),
    .CLK(clknet_leaf_30_user_clock2),
    .Q(\iram_latched[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3268_ (.D(_0049_),
    .CLK(clknet_leaf_31_user_clock2),
    .Q(\iram_latched[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3269_ (.D(_0050_),
    .CLK(clknet_leaf_31_user_clock2),
    .Q(\iram_latched[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3270_ (.D(_0051_),
    .CLK(clknet_leaf_31_user_clock2),
    .Q(\iram_latched[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3271_ (.D(_0052_),
    .CLK(clknet_leaf_30_user_clock2),
    .Q(\iram_latched[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3272_ (.D(_0053_),
    .CLK(clknet_leaf_30_user_clock2),
    .Q(\iram_latched[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3273_ (.D(_0054_),
    .CLK(clknet_leaf_30_user_clock2),
    .Q(\iram_latched[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3274_ (.D(_0055_),
    .CLK(clknet_leaf_29_user_clock2),
    .Q(\iram_latched[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3275_ (.D(_0056_),
    .CLK(clknet_leaf_29_user_clock2),
    .Q(\iram_latched[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3276_ (.D(_0057_),
    .CLK(clknet_leaf_29_user_clock2),
    .Q(\iram_latched[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3277_ (.D(_0058_),
    .CLK(clknet_leaf_28_user_clock2),
    .Q(\iram_latched[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3278_ (.D(_0059_),
    .CLK(clknet_leaf_29_user_clock2),
    .Q(\iram_latched[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3279_ (.D(_0060_),
    .CLK(clknet_leaf_30_user_clock2),
    .Q(\iram_latched[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3280_ (.D(_0061_),
    .CLK(clknet_leaf_33_user_clock2),
    .Q(iram_wb_ack_del),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3281_ (.D(_0062_),
    .CLK(clknet_leaf_50_user_clock2),
    .Q(\clk_div.res_clk ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3282_ (.D(_0063_),
    .CLK(clknet_leaf_42_user_clock2),
    .Q(\clk_div.next_div_buff[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3283_ (.D(_0064_),
    .CLK(clknet_leaf_43_user_clock2),
    .Q(\clk_div.next_div_buff[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3284_ (.D(_0065_),
    .CLK(clknet_leaf_42_user_clock2),
    .Q(\clk_div.next_div_buff[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3285_ (.D(_0066_),
    .CLK(clknet_leaf_43_user_clock2),
    .Q(\clk_div.next_div_buff[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3286_ (.D(_0067_),
    .CLK(clknet_leaf_43_user_clock2),
    .Q(\clk_div.next_div_val ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3287_ (.D(_0068_),
    .CLK(clknet_leaf_41_user_clock2),
    .Q(\clk_div.curr_div[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3288_ (.D(_0069_),
    .CLK(clknet_leaf_43_user_clock2),
    .Q(\clk_div.curr_div[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3289_ (.D(_0070_),
    .CLK(clknet_leaf_42_user_clock2),
    .Q(\clk_div.curr_div[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3290_ (.D(_0071_),
    .CLK(clknet_leaf_43_user_clock2),
    .Q(\clk_div.curr_div[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3291_ (.D(net539),
    .CLK(clknet_leaf_50_user_clock2),
    .Q(\clk_div.clock_sel_r ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3292_ (.D(_0072_),
    .CLK(clknet_4_1_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3293_ (.D(_0073_),
    .CLK(clknet_4_1_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3294_ (.D(_0074_),
    .CLK(clknet_4_1_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3295_ (.D(_0075_),
    .CLK(clknet_4_3_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3296_ (.D(_0076_),
    .CLK(clknet_4_8_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3297_ (.D(_0077_),
    .CLK(clknet_4_8_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3298_ (.D(_0078_),
    .CLK(clknet_4_10_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3299_ (.D(_0079_),
    .CLK(clknet_4_10_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3300_ (.D(_0080_),
    .CLK(clknet_4_10_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3301_ (.D(_0081_),
    .CLK(clknet_4_10_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3302_ (.D(_0082_),
    .CLK(clknet_4_10_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3303_ (.D(_0083_),
    .CLK(clknet_4_10_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3304_ (.D(_0084_),
    .CLK(clknet_4_10_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3305_ (.D(_0085_),
    .CLK(clknet_4_11_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3306_ (.D(_0086_),
    .CLK(clknet_4_11_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3307_ (.D(_0087_),
    .CLK(clknet_4_11_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3308_ (.D(_0088_),
    .CLK(clknet_4_11_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[16] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3309_ (.D(_0089_),
    .CLK(clknet_4_11_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[17] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3310_ (.D(_0090_),
    .CLK(clknet_4_11_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[18] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3311_ (.D(_0091_),
    .CLK(clknet_4_14_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[19] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3312_ (.D(_0092_),
    .CLK(clknet_4_14_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[20] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3313_ (.D(_0093_),
    .CLK(clknet_4_12_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[21] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3314_ (.D(_0094_),
    .CLK(clknet_4_11_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[22] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3315_ (.D(_0095_),
    .CLK(clknet_4_8_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[23] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3316_ (.D(_0096_),
    .CLK(clknet_4_10_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[24] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3317_ (.D(_0097_),
    .CLK(clknet_4_10_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[25] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3318_ (.D(_0098_),
    .CLK(clknet_4_10_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[26] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3319_ (.D(_0099_),
    .CLK(clknet_4_8_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[27] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3320_ (.D(_0100_),
    .CLK(clknet_4_11_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[28] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3321_ (.D(_0101_),
    .CLK(clknet_4_9_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[29] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3322_ (.D(_0102_),
    .CLK(clknet_4_9_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[30] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3323_ (.D(_0103_),
    .CLK(clknet_4_8_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[31] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3324_ (.D(_0104_),
    .CLK(clknet_4_8_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[32] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3325_ (.D(_0105_),
    .CLK(clknet_4_8_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[33] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3326_ (.D(_0106_),
    .CLK(clknet_4_6_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[34] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3327_ (.D(_0107_),
    .CLK(clknet_4_6_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[35] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3328_ (.D(_0108_),
    .CLK(clknet_4_6_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[36] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3329_ (.D(_0109_),
    .CLK(clknet_4_7_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[37] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3330_ (.D(_0110_),
    .CLK(clknet_4_7_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[38] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3331_ (.D(_0111_),
    .CLK(clknet_4_6_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[39] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3332_ (.D(_0112_),
    .CLK(clknet_4_6_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[40] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3333_ (.D(_0113_),
    .CLK(clknet_4_6_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[41] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3334_ (.D(_0114_),
    .CLK(clknet_4_4_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[42] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3335_ (.D(_0115_),
    .CLK(clknet_4_4_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[43] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3336_ (.D(_0116_),
    .CLK(clknet_4_1_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[44] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3337_ (.D(_0117_),
    .CLK(clknet_4_4_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[45] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3338_ (.D(_0118_),
    .CLK(clknet_4_1_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_data[46] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3339_ (.D(_0119_),
    .CLK(clknet_leaf_5_user_clock2),
    .Q(\wb_cross_clk.prev_ack ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3340_ (.D(_0120_),
    .CLK(clknet_leaf_50_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_xfer_xor_flag ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3341_ (.D(_0121_),
    .CLK(clknet_4_0_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3342_ (.D(_0122_),
    .CLK(clknet_4_3_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3343_ (.D(_0123_),
    .CLK(clknet_4_8_0_net196),
    .Q(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3344_ (.D(_0124_),
    .CLK(clknet_leaf_32_user_clock2),
    .Q(\wb_cross_clk.msy_xor_ack ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3345_ (.D(_0125_),
    .CLK(clknet_leaf_21_user_clock2),
    .Q(\wb_cross_clk.msy_xor_err ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3346_ (.D(_0126_),
    .CLK(clknet_leaf_32_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3347_ (.D(_0127_),
    .CLK(clknet_leaf_29_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3348_ (.D(_0128_),
    .CLK(clknet_leaf_29_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3349_ (.D(_0129_),
    .CLK(clknet_leaf_30_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3350_ (.D(_0130_),
    .CLK(clknet_leaf_29_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3351_ (.D(_0131_),
    .CLK(clknet_leaf_26_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3352_ (.D(_0132_),
    .CLK(clknet_leaf_26_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3353_ (.D(_0133_),
    .CLK(clknet_leaf_26_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3354_ (.D(_0134_),
    .CLK(clknet_leaf_24_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3355_ (.D(_0135_),
    .CLK(clknet_leaf_24_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3356_ (.D(_0136_),
    .CLK(clknet_leaf_17_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3357_ (.D(_0137_),
    .CLK(clknet_leaf_17_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3358_ (.D(_0138_),
    .CLK(clknet_leaf_17_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3359_ (.D(_0139_),
    .CLK(clknet_leaf_17_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3360_ (.D(_0140_),
    .CLK(clknet_leaf_23_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3361_ (.D(_0141_),
    .CLK(clknet_leaf_23_user_clock2),
    .Q(\wb_cross_clk.m_wb_i_dat[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3362_ (.D(_0142_),
    .CLK(clknet_leaf_1_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3363_ (.D(_0143_),
    .CLK(clknet_leaf_1_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3364_ (.D(_0144_),
    .CLK(clknet_leaf_1_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3365_ (.D(_0145_),
    .CLK(clknet_leaf_45_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3366_ (.D(_0146_),
    .CLK(clknet_leaf_45_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3367_ (.D(_0147_),
    .CLK(clknet_leaf_42_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3368_ (.D(_0148_),
    .CLK(clknet_leaf_42_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3369_ (.D(_0149_),
    .CLK(clknet_leaf_39_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3370_ (.D(_0150_),
    .CLK(clknet_leaf_39_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3371_ (.D(_0151_),
    .CLK(clknet_leaf_40_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3372_ (.D(_0152_),
    .CLK(clknet_leaf_39_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3373_ (.D(_0153_),
    .CLK(clknet_leaf_38_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3374_ (.D(_0154_),
    .CLK(clknet_leaf_37_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3375_ (.D(_0155_),
    .CLK(clknet_leaf_37_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3376_ (.D(_0156_),
    .CLK(clknet_leaf_31_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3377_ (.D(_0157_),
    .CLK(clknet_leaf_31_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3378_ (.D(_0158_),
    .CLK(clknet_leaf_37_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[16] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3379_ (.D(_0159_),
    .CLK(clknet_leaf_37_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[17] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3380_ (.D(_0160_),
    .CLK(clknet_leaf_31_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[18] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3381_ (.D(_0161_),
    .CLK(clknet_leaf_31_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[19] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3382_ (.D(_0162_),
    .CLK(clknet_leaf_31_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[20] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3383_ (.D(_0163_),
    .CLK(clknet_leaf_31_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[21] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3384_ (.D(_0164_),
    .CLK(clknet_leaf_35_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[22] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3385_ (.D(_0165_),
    .CLK(clknet_leaf_38_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[23] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3386_ (.D(_0166_),
    .CLK(clknet_leaf_39_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[24] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3387_ (.D(_0167_),
    .CLK(clknet_leaf_38_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[25] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3388_ (.D(_0168_),
    .CLK(clknet_leaf_35_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[26] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3389_ (.D(_0169_),
    .CLK(clknet_leaf_45_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[27] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3390_ (.D(_0170_),
    .CLK(clknet_leaf_36_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[28] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3391_ (.D(_0171_),
    .CLK(clknet_leaf_36_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[29] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3392_ (.D(_0172_),
    .CLK(clknet_2_2__leaf_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[30] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3393_ (.D(_0173_),
    .CLK(clknet_leaf_33_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[31] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3394_ (.D(_0174_),
    .CLK(clknet_leaf_33_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[32] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3395_ (.D(_0175_),
    .CLK(clknet_leaf_45_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[33] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3396_ (.D(_0176_),
    .CLK(clknet_leaf_46_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[34] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3397_ (.D(_0177_),
    .CLK(clknet_leaf_46_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[35] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3398_ (.D(_0178_),
    .CLK(clknet_leaf_46_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[36] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3399_ (.D(_0179_),
    .CLK(clknet_leaf_46_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[37] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3400_ (.D(_0180_),
    .CLK(clknet_leaf_6_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[38] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3401_ (.D(_0181_),
    .CLK(clknet_leaf_47_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[39] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3402_ (.D(_0182_),
    .CLK(clknet_leaf_47_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[40] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3403_ (.D(_0183_),
    .CLK(clknet_2_0__leaf_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[41] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3404_ (.D(_0184_),
    .CLK(clknet_leaf_47_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[42] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3405_ (.D(_0185_),
    .CLK(clknet_leaf_5_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[43] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3406_ (.D(_0186_),
    .CLK(clknet_leaf_5_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[44] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3407_ (.D(_0187_),
    .CLK(clknet_leaf_47_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[45] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3408_ (.D(_0188_),
    .CLK(clknet_leaf_5_user_clock2),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[46] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3409_ (.D(_0189_),
    .CLK(clknet_4_1_0_net196),
    .Q(\wb_cross_clk.s_m_sync.s_xfer_xor_flag ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3410_ (.D(_0190_),
    .CLK(clknet_leaf_47_user_clock2),
    .Q(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3411_ (.D(_0191_),
    .CLK(clknet_leaf_21_user_clock2),
    .Q(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3412_ (.D(_0192_),
    .CLK(clknet_leaf_22_user_clock2),
    .Q(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3413_ (.D(_0193_),
    .CLK(clknet_leaf_5_user_clock2),
    .Q(\wb_cross_clk.prev_stb ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3414_ (.D(_0194_),
    .CLK(clknet_leaf_21_user_clock2),
    .Q(\wb_cross_clk.prev_xor_err ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3415_ (.D(_0195_),
    .CLK(clknet_leaf_0_user_clock2),
    .Q(\wb_cross_clk.m_new_req_flag ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3416_ (.D(_0196_),
    .CLK(clknet_leaf_1_user_clock2),
    .Q(\wb_cross_clk.m_burst_cnt[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3417_ (.D(_0197_),
    .CLK(clknet_leaf_2_user_clock2),
    .Q(\wb_cross_clk.m_burst_cnt[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3418_ (.D(_0198_),
    .CLK(clknet_leaf_1_user_clock2),
    .Q(\wb_cross_clk.m_burst_cnt[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3419_ (.D(_0199_),
    .CLK(clknet_leaf_0_user_clock2),
    .Q(\wb_cross_clk.m_burst_cnt[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3420_ (.D(_0200_),
    .CLK(clknet_4_0_0_net196),
    .Q(\wb_cross_clk.s_burst_cnt[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3421_ (.D(_0201_),
    .CLK(clknet_4_0_0_net196),
    .Q(\wb_cross_clk.s_burst_cnt[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3422_ (.D(_0202_),
    .CLK(clknet_4_1_0_net196),
    .Q(\wb_cross_clk.s_burst_cnt[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3423_ (.D(_0203_),
    .CLK(clknet_4_3_0_net196),
    .Q(\wb_cross_clk.s_burst_cnt[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3424_ (.D(_0204_),
    .CLK(clknet_4_1_0_net196),
    .Q(\wb_cross_clk.ack_next_hold ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3425_ (.D(_0205_),
    .CLK(clknet_4_3_0_net196),
    .Q(\wb_cross_clk.err_xor_flag ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3426_ (.D(_0206_),
    .CLK(clknet_4_14_0_net196),
    .Q(\wb_cross_clk.ack_xor_flag ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3427_ (.D(_0207_),
    .CLK(clknet_leaf_32_user_clock2),
    .Q(\wb_cross_clk.prev_xor_ack ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3428_ (.D(_0208_),
    .CLK(clknet_4_0_0_net196),
    .Q(\wb_cross_clk.prev_xor_newreq ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3429_ (.D(_0209_),
    .CLK(clknet_4_2_0_net196),
    .Q(\wb_compressor.l_we ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3430_ (.D(net489),
    .CLK(clknet_4_0_0_net196),
    .Q(\wb_compressor.burst_end[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3431_ (.D(_0211_),
    .CLK(clknet_4_0_0_net196),
    .Q(\wb_compressor.burst_end[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3432_ (.D(_0212_),
    .CLK(clknet_4_15_0_net196),
    .Q(\wb_compressor.wb_i_dat[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3433_ (.D(_0213_),
    .CLK(clknet_4_15_0_net196),
    .Q(\wb_compressor.wb_i_dat[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3434_ (.D(_0214_),
    .CLK(clknet_4_15_0_net196),
    .Q(\wb_compressor.wb_i_dat[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3435_ (.D(_0215_),
    .CLK(clknet_4_14_0_net196),
    .Q(\wb_compressor.wb_i_dat[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3436_ (.D(_0216_),
    .CLK(clknet_4_15_0_net196),
    .Q(\wb_compressor.wb_i_dat[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3437_ (.D(_0217_),
    .CLK(clknet_4_15_0_net196),
    .Q(\wb_compressor.wb_i_dat[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3438_ (.D(_0218_),
    .CLK(clknet_4_15_0_net196),
    .Q(\wb_compressor.wb_i_dat[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3439_ (.D(_0219_),
    .CLK(clknet_4_13_0_net196),
    .Q(\wb_compressor.wb_i_dat[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3440_ (.D(_0220_),
    .CLK(clknet_4_13_0_net196),
    .Q(\wb_compressor.wb_i_dat[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3441_ (.D(_0221_),
    .CLK(clknet_4_13_0_net196),
    .Q(\wb_compressor.wb_i_dat[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3442_ (.D(_0222_),
    .CLK(clknet_4_5_0_net196),
    .Q(\wb_compressor.wb_i_dat[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3443_ (.D(_0223_),
    .CLK(clknet_4_5_0_net196),
    .Q(\wb_compressor.wb_i_dat[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3444_ (.D(_0224_),
    .CLK(clknet_4_5_0_net196),
    .Q(\wb_compressor.wb_i_dat[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3445_ (.D(_0225_),
    .CLK(clknet_4_5_0_net196),
    .Q(\wb_compressor.wb_i_dat[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3446_ (.D(_0226_),
    .CLK(clknet_4_7_0_net196),
    .Q(\wb_compressor.wb_i_dat[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3447_ (.D(_0227_),
    .CLK(clknet_4_12_0_net196),
    .Q(\wb_compressor.wb_i_dat[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3448_ (.D(_0228_),
    .CLK(clknet_4_6_0_net196),
    .Q(\wb_compressor.wb_err ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3449_ (.D(_0229_),
    .CLK(clknet_4_6_0_net196),
    .Q(\wb_compressor.wb_ack ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3450_ (.D(_0230_),
    .CLK(clknet_leaf_0_user_clock2),
    .Q(\sspi.sy_clk[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3451_ (.D(_0231_),
    .CLK(clknet_leaf_0_user_clock2),
    .Q(\sspi.sy_clk[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3452_ (.D(_0232_),
    .CLK(clknet_leaf_0_user_clock2),
    .Q(\sspi.sy_clk[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3453_ (.D(_0233_),
    .CLK(clknet_leaf_0_user_clock2),
    .Q(\sspi.sy_clk[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3454_ (.D(_0234_),
    .CLK(clknet_4_3_0_net196),
    .Q(net168),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3455_ (.D(_0235_),
    .CLK(clknet_4_3_0_net196),
    .Q(net202),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3456_ (.D(_0236_),
    .CLK(clknet_4_9_0_net196),
    .Q(net176),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3457_ (.D(_0237_),
    .CLK(clknet_4_9_0_net196),
    .Q(net177),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3458_ (.D(_0238_),
    .CLK(clknet_4_14_0_net196),
    .Q(net178),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3459_ (.D(_0239_),
    .CLK(clknet_4_14_0_net196),
    .Q(net179),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3460_ (.D(_0240_),
    .CLK(clknet_4_14_0_net196),
    .Q(net180),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3461_ (.D(_0241_),
    .CLK(clknet_4_12_0_net196),
    .Q(net181),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3462_ (.D(_0242_),
    .CLK(clknet_4_9_0_net196),
    .Q(net182),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3463_ (.D(_0243_),
    .CLK(clknet_4_9_0_net196),
    .Q(net183),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3464_ (.D(_0244_),
    .CLK(clknet_4_14_0_net196),
    .Q(net184),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3465_ (.D(_0245_),
    .CLK(clknet_4_14_0_net196),
    .Q(net185),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3466_ (.D(_0246_),
    .CLK(clknet_4_12_0_net196),
    .Q(net187),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3467_ (.D(_0247_),
    .CLK(clknet_4_12_0_net196),
    .Q(net188),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3468_ (.D(_0248_),
    .CLK(clknet_4_12_0_net196),
    .Q(net189),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3469_ (.D(_0249_),
    .CLK(clknet_4_12_0_net196),
    .Q(net190),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3470_ (.D(_0250_),
    .CLK(clknet_4_12_0_net196),
    .Q(net191),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3471_ (.D(_0251_),
    .CLK(clknet_4_12_0_net196),
    .Q(net192),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3472_ (.D(_0010_),
    .CLK(clknet_4_2_0_net196),
    .Q(\wb_compressor.state[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3473_ (.D(_0000_),
    .CLK(clknet_4_2_0_net196),
    .Q(\wb_compressor.state[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3474_ (.D(_0011_),
    .CLK(clknet_4_3_0_net196),
    .Q(\wb_compressor.state[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3475_ (.D(_0001_),
    .CLK(clknet_4_3_0_net196),
    .Q(\wb_compressor.state[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3476_ (.D(_0012_),
    .CLK(clknet_4_2_0_net196),
    .Q(\wb_compressor.state[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3477_ (.D(_0013_),
    .CLK(clknet_4_2_0_net196),
    .Q(\wb_compressor.state[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _3478_ (.D(_0014_),
    .CLK(clknet_4_3_0_net196),
    .Q(\wb_compressor.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3479_ (.D(_0002_),
    .CLK(clknet_leaf_5_user_clock2),
    .Q(\sspi.state[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3480_ (.D(_0003_),
    .CLK(clknet_leaf_2_user_clock2),
    .Q(\sspi.state[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3481_ (.D(_0004_),
    .CLK(clknet_leaf_3_user_clock2),
    .Q(\sspi.state[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3482_ (.D(_0005_),
    .CLK(clknet_leaf_2_user_clock2),
    .Q(\sspi.state[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3483_ (.D(_0006_),
    .CLK(clknet_leaf_3_user_clock2),
    .Q(\sspi.state[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3484_ (.D(_0007_),
    .CLK(clknet_leaf_2_user_clock2),
    .Q(\sspi.state[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3485_ (.D(_0008_),
    .CLK(clknet_leaf_3_user_clock2),
    .Q(\sspi.state[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3486_ (.D(_0009_),
    .CLK(clknet_leaf_2_user_clock2),
    .Q(\sspi.state[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3487_ (.D(_0252_),
    .CLK(clknet_leaf_5_user_clock2),
    .Q(\sspi.resp_err ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _3488_ (.D(_0253_),
    .CLK(clknet_leaf_12_user_clock2),
    .Q(\sspi.bit_cnt[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _3489_ (.D(_0254_),
    .CLK(clknet_leaf_11_user_clock2),
    .Q(\sspi.bit_cnt[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3490_ (.D(_0255_),
    .CLK(clknet_leaf_12_user_clock2),
    .Q(\sspi.bit_cnt[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _3491_ (.D(_0256_),
    .CLK(clknet_leaf_10_user_clock2),
    .Q(\sspi.bit_cnt[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3492_ (.D(_0257_),
    .CLK(clknet_leaf_10_user_clock2),
    .Q(\sspi.bit_cnt[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3493_ (.D(_0258_),
    .CLK(clknet_leaf_18_user_clock2),
    .Q(\sspi.res_data[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3494_ (.D(_0259_),
    .CLK(clknet_leaf_23_user_clock2),
    .Q(\sspi.res_data[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3495_ (.D(_0260_),
    .CLK(clknet_leaf_23_user_clock2),
    .Q(\sspi.res_data[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3496_ (.D(_0261_),
    .CLK(clknet_leaf_23_user_clock2),
    .Q(\sspi.res_data[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3497_ (.D(_0262_),
    .CLK(clknet_leaf_22_user_clock2),
    .Q(\sspi.res_data[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3498_ (.D(_0263_),
    .CLK(clknet_leaf_26_user_clock2),
    .Q(\sspi.res_data[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3499_ (.D(_0264_),
    .CLK(clknet_leaf_23_user_clock2),
    .Q(\sspi.res_data[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3500_ (.D(_0265_),
    .CLK(clknet_leaf_16_user_clock2),
    .Q(\sspi.res_data[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3501_ (.D(_0266_),
    .CLK(clknet_leaf_16_user_clock2),
    .Q(\sspi.res_data[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3502_ (.D(_0267_),
    .CLK(clknet_leaf_16_user_clock2),
    .Q(\sspi.res_data[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3503_ (.D(_0268_),
    .CLK(clknet_leaf_17_user_clock2),
    .Q(\sspi.res_data[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3504_ (.D(_0269_),
    .CLK(clknet_leaf_18_user_clock2),
    .Q(\sspi.res_data[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3505_ (.D(_0270_),
    .CLK(clknet_leaf_17_user_clock2),
    .Q(\sspi.res_data[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3506_ (.D(_0271_),
    .CLK(clknet_leaf_18_user_clock2),
    .Q(\sspi.res_data[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3507_ (.D(_0272_),
    .CLK(clknet_leaf_18_user_clock2),
    .Q(\sspi.res_data[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3508_ (.D(_0273_),
    .CLK(clknet_leaf_18_user_clock2),
    .Q(\sspi.res_data[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3509_ (.D(_0274_),
    .CLK(clknet_leaf_13_user_clock2),
    .Q(\sspi.req_data[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3510_ (.D(_0275_),
    .CLK(clknet_leaf_12_user_clock2),
    .Q(\sspi.req_data[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3511_ (.D(_0276_),
    .CLK(clknet_leaf_12_user_clock2),
    .Q(\sspi.req_data[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3512_ (.D(_0277_),
    .CLK(clknet_leaf_13_user_clock2),
    .Q(\sspi.req_data[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3513_ (.D(_0278_),
    .CLK(clknet_leaf_12_user_clock2),
    .Q(\sspi.req_data[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3514_ (.D(_0279_),
    .CLK(clknet_leaf_16_user_clock2),
    .Q(\sspi.req_data[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3515_ (.D(_0280_),
    .CLK(clknet_leaf_16_user_clock2),
    .Q(\sspi.req_data[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3516_ (.D(_0281_),
    .CLK(clknet_leaf_10_user_clock2),
    .Q(\sspi.req_data[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3517_ (.D(_0282_),
    .CLK(clknet_leaf_16_user_clock2),
    .Q(\sspi.req_data[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3518_ (.D(_0283_),
    .CLK(clknet_leaf_8_user_clock2),
    .Q(\sspi.req_data[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3519_ (.D(_0284_),
    .CLK(clknet_leaf_18_user_clock2),
    .Q(\sspi.req_data[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3520_ (.D(_0285_),
    .CLK(clknet_leaf_19_user_clock2),
    .Q(\sspi.req_data[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3521_ (.D(_0286_),
    .CLK(clknet_leaf_19_user_clock2),
    .Q(\sspi.req_data[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3522_ (.D(_0287_),
    .CLK(clknet_leaf_16_user_clock2),
    .Q(\sspi.req_data[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3523_ (.D(_0288_),
    .CLK(clknet_leaf_16_user_clock2),
    .Q(\sspi.req_data[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3524_ (.D(_0289_),
    .CLK(clknet_leaf_12_user_clock2),
    .Q(\sspi.req_data[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3525_ (.D(_0290_),
    .CLK(clknet_leaf_9_user_clock2),
    .Q(\sspi.req_addr[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3526_ (.D(_0291_),
    .CLK(clknet_leaf_9_user_clock2),
    .Q(\sspi.req_addr[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3527_ (.D(_0292_),
    .CLK(clknet_leaf_9_user_clock2),
    .Q(\sspi.req_addr[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3528_ (.D(_0293_),
    .CLK(clknet_leaf_8_user_clock2),
    .Q(\sspi.req_addr[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3529_ (.D(_0294_),
    .CLK(clknet_leaf_9_user_clock2),
    .Q(\sspi.req_addr[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3530_ (.D(_0295_),
    .CLK(clknet_leaf_7_user_clock2),
    .Q(\sspi.req_addr[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3531_ (.D(_0296_),
    .CLK(clknet_leaf_8_user_clock2),
    .Q(\sspi.req_addr[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3532_ (.D(_0297_),
    .CLK(clknet_leaf_11_user_clock2),
    .Q(\sspi.req_addr[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3533_ (.D(_0298_),
    .CLK(clknet_leaf_8_user_clock2),
    .Q(\sspi.req_addr[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3534_ (.D(_0299_),
    .CLK(clknet_leaf_8_user_clock2),
    .Q(\sspi.req_addr[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3535_ (.D(_0300_),
    .CLK(clknet_leaf_19_user_clock2),
    .Q(\sspi.req_addr[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3536_ (.D(_0301_),
    .CLK(clknet_leaf_19_user_clock2),
    .Q(\sspi.req_addr[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3537_ (.D(_0302_),
    .CLK(clknet_leaf_19_user_clock2),
    .Q(\sspi.req_addr[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3538_ (.D(_0303_),
    .CLK(clknet_leaf_8_user_clock2),
    .Q(\sspi.req_addr[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3539_ (.D(_0304_),
    .CLK(clknet_leaf_11_user_clock2),
    .Q(\sspi.req_addr[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3540_ (.D(_0305_),
    .CLK(clknet_leaf_9_user_clock2),
    .Q(\sspi.req_addr[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3541_ (.D(_0306_),
    .CLK(clknet_leaf_9_user_clock2),
    .Q(\sspi.req_addr[16] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3542_ (.D(_0307_),
    .CLK(clknet_leaf_8_user_clock2),
    .Q(\sspi.req_addr[17] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3543_ (.D(_0308_),
    .CLK(clknet_leaf_4_user_clock2),
    .Q(\sspi.req_addr[18] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3544_ (.D(_0309_),
    .CLK(clknet_leaf_7_user_clock2),
    .Q(\sspi.req_addr[19] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3545_ (.D(_0310_),
    .CLK(clknet_leaf_4_user_clock2),
    .Q(\sspi.req_addr[20] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3546_ (.D(_0311_),
    .CLK(clknet_leaf_7_user_clock2),
    .Q(\sspi.req_addr[21] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3547_ (.D(_0312_),
    .CLK(clknet_leaf_8_user_clock2),
    .Q(\sspi.req_addr[22] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3548_ (.D(_0313_),
    .CLK(clknet_leaf_9_user_clock2),
    .Q(\sspi.req_addr[23] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3549_ (.D(_0314_),
    .CLK(clknet_leaf_6_user_clock2),
    .Q(\m_arbiter.wb0_we ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3550_ (.D(_0315_),
    .CLK(clknet_leaf_14_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3551_ (.D(_0316_),
    .CLK(clknet_leaf_13_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3552_ (.D(_0317_),
    .CLK(clknet_leaf_13_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3553_ (.D(_0318_),
    .CLK(clknet_leaf_14_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3554_ (.D(_0319_),
    .CLK(clknet_leaf_13_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3555_ (.D(_0320_),
    .CLK(clknet_leaf_15_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3556_ (.D(_0321_),
    .CLK(clknet_leaf_14_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3557_ (.D(_0322_),
    .CLK(clknet_leaf_13_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3558_ (.D(_0323_),
    .CLK(clknet_leaf_16_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3559_ (.D(_0324_),
    .CLK(clknet_leaf_21_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3560_ (.D(_0325_),
    .CLK(clknet_leaf_18_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3561_ (.D(_0326_),
    .CLK(clknet_leaf_18_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3562_ (.D(_0327_),
    .CLK(clknet_leaf_23_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3563_ (.D(_0328_),
    .CLK(clknet_leaf_15_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3564_ (.D(_0329_),
    .CLK(clknet_leaf_15_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3565_ (.D(_0330_),
    .CLK(clknet_leaf_14_user_clock2),
    .Q(\m_arbiter.wb0_o_dat[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3566_ (.D(_0331_),
    .CLK(clknet_leaf_41_user_clock2),
    .Q(\clk_div.cnt[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3567_ (.D(_0332_),
    .CLK(clknet_leaf_41_user_clock2),
    .Q(\clk_div.cnt[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3568_ (.D(_0333_),
    .CLK(clknet_leaf_41_user_clock2),
    .Q(\clk_div.cnt[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3569_ (.D(_0334_),
    .CLK(clknet_leaf_41_user_clock2),
    .Q(\clk_div.cnt[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3570_ (.D(_0335_),
    .CLK(clknet_leaf_43_user_clock2),
    .Q(\clk_div.cnt[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3571_ (.D(_0336_),
    .CLK(clknet_leaf_41_user_clock2),
    .Q(\clk_div.cnt[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3572_ (.D(_0337_),
    .CLK(clknet_leaf_41_user_clock2),
    .Q(\clk_div.cnt[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3573_ (.D(_0338_),
    .CLK(clknet_leaf_44_user_clock2),
    .Q(\clk_div.cnt[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3574_ (.D(_0339_),
    .CLK(clknet_leaf_44_user_clock2),
    .Q(\clk_div.cnt[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3575_ (.D(_0340_),
    .CLK(clknet_leaf_44_user_clock2),
    .Q(\clk_div.cnt[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3576_ (.D(_0341_),
    .CLK(clknet_leaf_44_user_clock2),
    .Q(\clk_div.cnt[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3577_ (.D(_0342_),
    .CLK(clknet_leaf_44_user_clock2),
    .Q(\clk_div.cnt[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3578_ (.D(_0343_),
    .CLK(clknet_leaf_49_user_clock2),
    .Q(\clk_div.cnt[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3579_ (.D(_0344_),
    .CLK(clknet_leaf_49_user_clock2),
    .Q(\clk_div.cnt[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3580_ (.D(_0345_),
    .CLK(clknet_leaf_49_user_clock2),
    .Q(\clk_div.cnt[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3581_ (.D(_0346_),
    .CLK(clknet_leaf_49_user_clock2),
    .Q(\clk_div.cnt[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3582_ (.D(_0347_),
    .CLK(clknet_leaf_5_user_clock2),
    .Q(\m_arbiter.i_wb0_cyc ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3583_ (.D(_0348_),
    .CLK(clknet_leaf_2_user_clock2),
    .Q(net195),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3584_ (.D(_0349_),
    .CLK(clknet_leaf_7_user_clock2),
    .Q(\m_arbiter.wb0_adr[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3585_ (.D(_0350_),
    .CLK(clknet_leaf_9_user_clock2),
    .Q(\m_arbiter.wb0_adr[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3586_ (.D(_0351_),
    .CLK(clknet_leaf_4_user_clock2),
    .Q(\m_arbiter.wb0_adr[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3587_ (.D(_0352_),
    .CLK(clknet_leaf_8_user_clock2),
    .Q(\m_arbiter.wb0_adr[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3588_ (.D(_0353_),
    .CLK(clknet_leaf_3_user_clock2),
    .Q(\m_arbiter.wb0_adr[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3589_ (.D(_0354_),
    .CLK(clknet_leaf_20_user_clock2),
    .Q(\m_arbiter.wb0_adr[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3590_ (.D(_0355_),
    .CLK(clknet_leaf_7_user_clock2),
    .Q(\m_arbiter.wb0_adr[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3591_ (.D(_0356_),
    .CLK(clknet_leaf_21_user_clock2),
    .Q(\m_arbiter.wb0_adr[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3592_ (.D(_0357_),
    .CLK(clknet_leaf_20_user_clock2),
    .Q(\m_arbiter.wb0_adr[8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3593_ (.D(_0358_),
    .CLK(clknet_leaf_7_user_clock2),
    .Q(\m_arbiter.wb0_adr[9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3594_ (.D(_0359_),
    .CLK(clknet_leaf_20_user_clock2),
    .Q(\m_arbiter.wb0_adr[10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3595_ (.D(_0360_),
    .CLK(clknet_leaf_19_user_clock2),
    .Q(\m_arbiter.wb0_adr[11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3596_ (.D(_0361_),
    .CLK(clknet_leaf_7_user_clock2),
    .Q(\m_arbiter.wb0_adr[12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3597_ (.D(_0362_),
    .CLK(clknet_leaf_20_user_clock2),
    .Q(\m_arbiter.wb0_adr[13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3598_ (.D(_0363_),
    .CLK(clknet_leaf_20_user_clock2),
    .Q(\m_arbiter.wb0_adr[14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3599_ (.D(_0364_),
    .CLK(clknet_leaf_20_user_clock2),
    .Q(\m_arbiter.wb0_adr[15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3600_ (.D(_0365_),
    .CLK(clknet_leaf_6_user_clock2),
    .Q(\m_arbiter.wb0_adr[16] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3601_ (.D(_0366_),
    .CLK(clknet_leaf_6_user_clock2),
    .Q(\m_arbiter.wb0_adr[17] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3602_ (.D(_0367_),
    .CLK(clknet_leaf_4_user_clock2),
    .Q(\m_arbiter.wb0_adr[18] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3603_ (.D(_0368_),
    .CLK(clknet_leaf_5_user_clock2),
    .Q(\m_arbiter.wb0_adr[19] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3604_ (.D(_0369_),
    .CLK(clknet_leaf_4_user_clock2),
    .Q(\m_arbiter.wb0_adr[20] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3605_ (.D(_0370_),
    .CLK(clknet_leaf_6_user_clock2),
    .Q(\m_arbiter.wb0_adr[21] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3606_ (.D(_0371_),
    .CLK(clknet_leaf_7_user_clock2),
    .Q(\m_arbiter.wb0_adr[22] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3607_ (.D(_0372_),
    .CLK(clknet_leaf_6_user_clock2),
    .Q(\m_arbiter.wb0_adr[23] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3608_ (.D(_0373_),
    .CLK(clknet_leaf_28_user_clock2),
    .Q(net151),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3609_ (.D(_0374_),
    .CLK(clknet_leaf_28_user_clock2),
    .Q(net162),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3610_ (.D(_0375_),
    .CLK(clknet_leaf_27_user_clock2),
    .Q(net169),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3611_ (.D(_0376_),
    .CLK(clknet_leaf_28_user_clock2),
    .Q(net170),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3612_ (.D(_0377_),
    .CLK(clknet_leaf_27_user_clock2),
    .Q(net171),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3613_ (.D(_0378_),
    .CLK(clknet_leaf_27_user_clock2),
    .Q(net172),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3614_ (.D(_0379_),
    .CLK(clknet_leaf_25_user_clock2),
    .Q(net173),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3615_ (.D(_0380_),
    .CLK(clknet_leaf_25_user_clock2),
    .Q(net174),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3616_ (.D(_0381_),
    .CLK(clknet_leaf_28_user_clock2),
    .Q(net175),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3617_ (.D(_0382_),
    .CLK(clknet_leaf_28_user_clock2),
    .Q(net186),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3618_ (.D(_0383_),
    .CLK(clknet_leaf_29_user_clock2),
    .Q(net194),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3619_ (.D(_0384_),
    .CLK(clknet_leaf_27_user_clock2),
    .Q(net197),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3620_ (.D(_0385_),
    .CLK(clknet_leaf_27_user_clock2),
    .Q(net198),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3621_ (.D(_0386_),
    .CLK(clknet_leaf_27_user_clock2),
    .Q(net199),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3622_ (.D(_0387_),
    .CLK(clknet_leaf_27_user_clock2),
    .Q(net200),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3623_ (.D(_0388_),
    .CLK(clknet_leaf_27_user_clock2),
    .Q(net201),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _3624_ (.D(net263),
    .SETN(_0015_),
    .CLK(clknet_leaf_50_user_clock2),
    .Q(\rst_soc_sync.reset_sync_ff[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3624__263 (.ZN(net263),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _3625_ (.D(\rst_soc_sync.reset_sync_ff[0] ),
    .SETN(_0016_),
    .CLK(clknet_leaf_50_user_clock2),
    .Q(\rst_soc_sync.reset_sync_ff[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _3626_ (.D(\rst_soc_sync.reset_sync_ff[1] ),
    .SETN(_0017_),
    .CLK(clknet_leaf_50_user_clock2),
    .Q(\rst_soc_sync.reset_sync_ff[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _3627_ (.D(\rst_soc_sync.reset_sync_ff[2] ),
    .SETN(_0018_),
    .CLK(clknet_leaf_50_user_clock2),
    .Q(net108),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _3628_ (.D(net264),
    .SETN(_0019_),
    .CLK(clknet_4_0_0_net196),
    .Q(\rst_cw_sync.reset_sync_ff[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3628__264 (.ZN(net264),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _3629_ (.D(\rst_cw_sync.reset_sync_ff[0] ),
    .SETN(_0020_),
    .CLK(clknet_4_0_0_net196),
    .Q(\rst_cw_sync.reset_sync_ff[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _3630_ (.D(\rst_cw_sync.reset_sync_ff[1] ),
    .SETN(_0021_),
    .CLK(clknet_4_0_0_net196),
    .Q(\rst_cw_sync.reset_sync_ff[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _3631_ (.D(\rst_cw_sync.reset_sync_ff[2] ),
    .SETN(_0022_),
    .CLK(clknet_4_0_0_net196),
    .Q(net193),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3632_ (.D(_0389_),
    .CLK(clknet_leaf_4_user_clock2),
    .Q(\m_arbiter.o_sel_sig ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3758_ (.I(clknet_leaf_13_user_clock2),
    .Z(net99),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3759_ (.I(clknet_leaf_24_user_clock2),
    .Z(net100),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3760_ (.I(clknet_leaf_24_user_clock2),
    .Z(net101),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3761_ (.I(clknet_leaf_13_user_clock2),
    .Z(net102),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3762_ (.I(clknet_leaf_24_user_clock2),
    .Z(net103),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3763_ (.I(clknet_leaf_13_user_clock2),
    .Z(net104),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3764_ (.I(clknet_leaf_40_user_clock2),
    .Z(net133),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3765_ (.I(net249),
    .Z(net152),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3766_ (.I(net249),
    .Z(net153),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3767_ (.I(net249),
    .Z(net154),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3768_ (.I(net249),
    .Z(net155),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3769_ (.I(net249),
    .Z(net156),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3770_ (.I(net249),
    .Z(net157),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3771_ (.I(net249),
    .Z(net158),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3772_ (.I(net249),
    .Z(net159),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3773_ (.I(net249),
    .Z(net160),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3774_ (.I(net249),
    .Z(net161),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3775_ (.I(net250),
    .Z(net163),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3776_ (.I(net250),
    .Z(net164),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3777_ (.I(net250),
    .Z(net165),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3778_ (.I(net250),
    .Z(net166),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3779_ (.I(net250),
    .Z(net167),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3780_ (.I(net250),
    .Z(net203),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_net196 (.I(net196),
    .Z(clknet_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_user_clock2 (.I(user_clock2),
    .Z(clknet_0_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_user_clock2 (.I(clknet_0_user_clock2),
    .Z(clknet_2_0__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_user_clock2 (.I(clknet_0_user_clock2),
    .Z(clknet_2_1__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_user_clock2 (.I(clknet_0_user_clock2),
    .Z(clknet_2_2__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_user_clock2 (.I(clknet_0_user_clock2),
    .Z(clknet_2_3__leaf_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_0_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_0_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_10_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_10_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_11_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_11_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_12_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_12_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_13_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_13_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_14_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_14_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_15_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_15_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_1_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_1_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_2_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_2_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_3_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_3_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_4_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_4_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_5_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_5_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_6_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_6_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_7_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_7_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_8_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_8_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_9_0_net196 (.I(clknet_0_net196),
    .Z(clknet_4_9_0_net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_user_clock2 (.I(clknet_2_0__leaf_user_clock2),
    .Z(clknet_leaf_0_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_10_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_11_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_12_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_13_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_14_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_15_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_16_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_17_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_18_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_19_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_user_clock2 (.I(clknet_2_0__leaf_user_clock2),
    .Z(clknet_leaf_1_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_20_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_user_clock2 (.I(clknet_2_3__leaf_user_clock2),
    .Z(clknet_leaf_21_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_user_clock2 (.I(clknet_2_3__leaf_user_clock2),
    .Z(clknet_leaf_22_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_user_clock2 (.I(clknet_2_3__leaf_user_clock2),
    .Z(clknet_leaf_23_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_user_clock2 (.I(clknet_2_3__leaf_user_clock2),
    .Z(clknet_leaf_24_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_user_clock2 (.I(clknet_2_3__leaf_user_clock2),
    .Z(clknet_leaf_25_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_user_clock2 (.I(clknet_2_3__leaf_user_clock2),
    .Z(clknet_leaf_26_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_user_clock2 (.I(clknet_2_3__leaf_user_clock2),
    .Z(clknet_leaf_27_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_user_clock2 (.I(clknet_2_3__leaf_user_clock2),
    .Z(clknet_leaf_28_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_user_clock2 (.I(clknet_2_3__leaf_user_clock2),
    .Z(clknet_leaf_29_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_user_clock2 (.I(clknet_2_0__leaf_user_clock2),
    .Z(clknet_leaf_2_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_user_clock2 (.I(clknet_2_3__leaf_user_clock2),
    .Z(clknet_leaf_30_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_user_clock2 (.I(clknet_2_3__leaf_user_clock2),
    .Z(clknet_leaf_31_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_user_clock2 (.I(clknet_2_3__leaf_user_clock2),
    .Z(clknet_leaf_32_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_user_clock2 (.I(clknet_2_2__leaf_user_clock2),
    .Z(clknet_leaf_33_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_user_clock2 (.I(clknet_2_2__leaf_user_clock2),
    .Z(clknet_leaf_35_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_user_clock2 (.I(clknet_2_2__leaf_user_clock2),
    .Z(clknet_leaf_36_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_user_clock2 (.I(clknet_2_2__leaf_user_clock2),
    .Z(clknet_leaf_37_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_user_clock2 (.I(clknet_2_2__leaf_user_clock2),
    .Z(clknet_leaf_38_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_user_clock2 (.I(clknet_2_2__leaf_user_clock2),
    .Z(clknet_leaf_39_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_user_clock2 (.I(clknet_2_0__leaf_user_clock2),
    .Z(clknet_leaf_3_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_user_clock2 (.I(clknet_2_2__leaf_user_clock2),
    .Z(clknet_leaf_40_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_user_clock2 (.I(clknet_2_2__leaf_user_clock2),
    .Z(clknet_leaf_41_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_user_clock2 (.I(clknet_2_2__leaf_user_clock2),
    .Z(clknet_leaf_42_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_user_clock2 (.I(clknet_2_2__leaf_user_clock2),
    .Z(clknet_leaf_43_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_user_clock2 (.I(clknet_2_2__leaf_user_clock2),
    .Z(clknet_leaf_44_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_user_clock2 (.I(clknet_2_2__leaf_user_clock2),
    .Z(clknet_leaf_45_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_user_clock2 (.I(clknet_2_2__leaf_user_clock2),
    .Z(clknet_leaf_46_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_user_clock2 (.I(clknet_2_0__leaf_user_clock2),
    .Z(clknet_leaf_47_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_user_clock2 (.I(clknet_2_0__leaf_user_clock2),
    .Z(clknet_leaf_49_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_user_clock2 (.I(clknet_2_0__leaf_user_clock2),
    .Z(clknet_leaf_4_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_user_clock2 (.I(clknet_2_0__leaf_user_clock2),
    .Z(clknet_leaf_50_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_user_clock2 (.I(clknet_2_0__leaf_user_clock2),
    .Z(clknet_leaf_5_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_user_clock2 (.I(clknet_2_0__leaf_user_clock2),
    .Z(clknet_leaf_6_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_7_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_8_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_user_clock2 (.I(clknet_2_1__leaf_user_clock2),
    .Z(clknet_leaf_9_user_clock2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout249 (.I(net250),
    .Z(net249),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout250 (.I(net168),
    .Z(net250),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold10 (.I(_0843_),
    .Z(net397),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold100 (.I(_1032_),
    .Z(net487),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold101 (.I(_1036_),
    .Z(net488),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold102 (.I(_0210_),
    .Z(net489),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold103 (.I(net526),
    .Z(net490),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold104 (.I(_0530_),
    .Z(net491),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold105 (.I(net108),
    .Z(net503),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold106 (.I(_1563_),
    .Z(net493),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold107 (.I(_1132_),
    .Z(net494),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold108 (.I(net538),
    .Z(net506),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold109 (.I(_1570_),
    .Z(net496),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold11 (.I(\wb_cross_clk.m_s_sync.s_data_ff[26] ),
    .Z(net398),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold110 (.I(_1163_),
    .Z(net497),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold111 (.I(_1164_),
    .Z(net498),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold112 (.I(\m_arbiter.wb0_we ),
    .Z(net499),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold113 (.I(net107),
    .Z(net508),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold114 (.I(_0396_),
    .Z(net501),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold115 (.I(_1138_),
    .Z(net502),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold116 (.I(net536),
    .Z(net511),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold117 (.I(_1564_),
    .Z(net504),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold118 (.I(_1127_),
    .Z(net505),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold119 (.I(\wb_cross_clk.m_s_sync.s_data_ff[0] ),
    .Z(net514),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold12 (.I(_0834_),
    .Z(net399),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold120 (.I(_1567_),
    .Z(net507),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold121 (.I(\wb_cross_clk.m_s_sync.s_data_ff[19] ),
    .Z(net517),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold122 (.I(_1582_),
    .Z(net509),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold123 (.I(_1150_),
    .Z(net510),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold124 (.I(\wb_cross_clk.m_s_sync.s_data_ff[21] ),
    .Z(net520),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold125 (.I(_1558_),
    .Z(net512),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold126 (.I(_1144_),
    .Z(net513),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold127 (.I(\wb_cross_clk.m_s_sync.s_data_ff[20] ),
    .Z(net523),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold128 (.I(_1581_),
    .Z(net515),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold129 (.I(_1156_),
    .Z(net516),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(\wb_cross_clk.m_s_sync.s_xfer_xor_flag ),
    .Z(net400),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold130 (.I(\clk_div.clock_sel ),
    .Z(net526),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold131 (.I(_1560_),
    .Z(net518),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold132 (.I(_1172_),
    .Z(net519),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold133 (.I(\wb_cross_clk.m_s_sync.s_data_ff[41] ),
    .Z(net527),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold134 (.I(_1572_),
    .Z(net521),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold135 (.I(_1168_),
    .Z(net522),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold136 (.I(\wb_cross_clk.m_s_sync.s_data_ff[30] ),
    .Z(net533),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold137 (.I(_1561_),
    .Z(net524),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold138 (.I(_1176_),
    .Z(net525),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold14 (.I(_0879_),
    .Z(net401),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold141 (.I(net130),
    .Z(net528),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold142 (.I(\embed_s_ff[0] ),
    .Z(net529),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold143 (.I(\disable_s_ff[0] ),
    .Z(net530),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold144 (.I(\m_arbiter.wb0_o_dat[0] ),
    .Z(net531),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold145 (.I(\split_s_ff[0] ),
    .Z(net532),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold147 (.I(net129),
    .Z(net534),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold148 (.I(\irq_s_ff[0] ),
    .Z(net535),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold149 (.I(net508),
    .Z(net536),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(\wb_cross_clk.m_s_sync.s_data_ff[40] ),
    .Z(net402),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold150 (.I(net390),
    .Z(net537),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold151 (.I(net503),
    .Z(net538),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold152 (.I(\clk_div.clock_sel ),
    .Z(net539),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(_0865_),
    .Z(net403),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(\wb_cross_clk.m_s_sync.s_data_ff[9] ),
    .Z(net404),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold18 (.I(_0796_),
    .Z(net405),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(\wb_cross_clk.m_s_sync.s_data_ff[39] ),
    .Z(net406),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(_0862_),
    .Z(net407),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(\wb_cross_clk.m_s_sync.s_data_ff[14] ),
    .Z(net408),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(_0808_),
    .Z(net409),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(\wb_cross_clk.m_s_sync.s_data_ff[25] ),
    .Z(net410),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(_0832_),
    .Z(net411),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(\wb_cross_clk.m_s_sync.s_data_ff[1] ),
    .Z(net412),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(_0778_),
    .Z(net413),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(\wb_cross_clk.m_s_sync.s_data_ff[11] ),
    .Z(net414),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(_0801_),
    .Z(net415),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(\wb_cross_clk.m_s_sync.s_data_ff[7] ),
    .Z(net416),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold3 (.I(net511),
    .Z(net390),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold30 (.I(_0791_),
    .Z(net417),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(\wb_cross_clk.m_s_sync.s_data_ff[8] ),
    .Z(net418),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(_0793_),
    .Z(net419),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(\wb_cross_clk.m_s_sync.s_data_ff[28] ),
    .Z(net420),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(_0839_),
    .Z(net421),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(\wb_cross_clk.m_s_sync.s_data_ff[22] ),
    .Z(net422),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(_0825_),
    .Z(net423),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(\wb_cross_clk.m_s_sync.s_data_ff[18] ),
    .Z(net424),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(_0816_),
    .Z(net425),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(\wb_cross_clk.m_s_sync.s_data_ff[3] ),
    .Z(net426),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 hold4 (.I(net391),
    .Z(inner_ext_irq),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(_0782_),
    .Z(net427),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(\wb_cross_clk.m_s_sync.s_data_ff[10] ),
    .Z(net428),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(_0798_),
    .Z(net429),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(\wb_cross_clk.m_s_sync.s_data_ff[23] ),
    .Z(net430),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(_0827_),
    .Z(net431),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(\wb_cross_clk.m_s_sync.s_data_ff[6] ),
    .Z(net432),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold46 (.I(_0789_),
    .Z(net433),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(\wb_cross_clk.m_s_sync.s_data_ff[15] ),
    .Z(net434),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold48 (.I(_0810_),
    .Z(net435),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(\wb_cross_clk.m_s_sync.s_data_ff[34] ),
    .Z(net436),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold5 (.I(net506),
    .Z(net392),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold50 (.I(_0853_),
    .Z(net437),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(\wb_cross_clk.m_s_sync.s_data_ff[35] ),
    .Z(net438),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold52 (.I(_0855_),
    .Z(net439),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(\wb_cross_clk.m_s_sync.s_data_ff[24] ),
    .Z(net440),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold54 (.I(_0830_),
    .Z(net441),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(\wb_cross_clk.m_s_sync.s_data_ff[4] ),
    .Z(net442),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold56 (.I(_0785_),
    .Z(net443),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(\wb_cross_clk.m_s_sync.s_data_ff[5] ),
    .Z(net444),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(_0787_),
    .Z(net445),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(\wb_cross_clk.m_s_sync.s_data_ff[36] ),
    .Z(net446),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 hold6 (.I(net393),
    .Z(inner_reset),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(_0857_),
    .Z(net447),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(\wb_cross_clk.m_s_sync.s_data_ff[33] ),
    .Z(net448),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold62 (.I(_0850_),
    .Z(net449),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(\wb_cross_clk.m_s_sync.s_data_ff[13] ),
    .Z(net450),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(_0805_),
    .Z(net451),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(\wb_cross_clk.m_s_sync.s_data_ff[12] ),
    .Z(net452),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold66 (.I(_0803_),
    .Z(net453),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(\wb_cross_clk.m_s_sync.s_data_ff[17] ),
    .Z(net454),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold68 (.I(_0814_),
    .Z(net455),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold69 (.I(\wb_cross_clk.m_s_sync.s_data_ff[31] ),
    .Z(net456),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold7 (.I(net527),
    .Z(net394),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(_0845_),
    .Z(net457),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(\wb_cross_clk.m_s_sync.s_data_ff[46] ),
    .Z(net458),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(_0877_),
    .Z(net459),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold73 (.I(\wb_cross_clk.m_s_sync.s_data_ff[42] ),
    .Z(net460),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold74 (.I(_0868_),
    .Z(net461),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold75 (.I(\wb_cross_clk.m_s_sync.s_data_ff[27] ),
    .Z(net462),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold76 (.I(_0837_),
    .Z(net463),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(\wb_cross_clk.m_s_sync.s_data_ff[32] ),
    .Z(net464),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold78 (.I(_0848_),
    .Z(net465),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold79 (.I(\wb_cross_clk.m_s_sync.s_data_ff[38] ),
    .Z(net466),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold8 (.I(_0866_),
    .Z(net395),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold80 (.I(_0860_),
    .Z(net467),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold81 (.I(\wb_cross_clk.m_s_sync.s_data_ff[44] ),
    .Z(net468),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(_0873_),
    .Z(net469),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold83 (.I(\wb_cross_clk.m_s_sync.s_data_ff[45] ),
    .Z(net470),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold84 (.I(_0875_),
    .Z(net471),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold85 (.I(\wb_cross_clk.m_s_sync.s_data_ff[29] ),
    .Z(net472),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold86 (.I(_0841_),
    .Z(net473),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold87 (.I(\wb_cross_clk.m_s_sync.s_data_ff[16] ),
    .Z(net474),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold88 (.I(_0812_),
    .Z(net475),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold89 (.I(\wb_cross_clk.m_s_sync.s_data_ff[37] ),
    .Z(net476),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold9 (.I(net533),
    .Z(net396),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold90 (.I(_0859_),
    .Z(net477),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold91 (.I(\wb_cross_clk.m_s_sync.s_data_ff[43] ),
    .Z(net478),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold92 (.I(_0871_),
    .Z(net479),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold93 (.I(\wb_cross_clk.m_s_sync.s_data_ff[2] ),
    .Z(net480),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold94 (.I(_0779_),
    .Z(net481),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold95 (.I(net514),
    .Z(net482),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold96 (.I(net517),
    .Z(net483),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold97 (.I(net523),
    .Z(net484),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold98 (.I(net520),
    .Z(net485),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold99 (.I(inner_wb_8_burst),
    .Z(net486),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1 (.I(inner_wb_4_burst),
    .Z(net1),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(inner_wb_adr[16]),
    .Z(net10),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(inner_wb_adr[17]),
    .Z(net11),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(inner_wb_adr[18]),
    .Z(net12),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(inner_wb_adr[19]),
    .Z(net13),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(inner_wb_adr[1]),
    .Z(net14),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(inner_wb_adr[20]),
    .Z(net15),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input16 (.I(inner_wb_adr[21]),
    .Z(net16),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(inner_wb_adr[22]),
    .Z(net17),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input18 (.I(inner_wb_adr[23]),
    .Z(net18),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(inner_wb_adr[2]),
    .Z(net19),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(net486),
    .Z(net2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(inner_wb_adr[3]),
    .Z(net20),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(inner_wb_adr[4]),
    .Z(net21),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input22 (.I(inner_wb_adr[5]),
    .Z(net22),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(inner_wb_adr[6]),
    .Z(net23),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input24 (.I(inner_wb_adr[7]),
    .Z(net24),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input25 (.I(inner_wb_adr[8]),
    .Z(net25),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(inner_wb_adr[9]),
    .Z(net26),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input27 (.I(inner_wb_cyc),
    .Z(net27),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(inner_wb_o_dat[0]),
    .Z(net28),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(inner_wb_o_dat[10]),
    .Z(net29),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input3 (.I(inner_wb_adr[0]),
    .Z(net3),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(inner_wb_o_dat[11]),
    .Z(net30),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(inner_wb_o_dat[12]),
    .Z(net31),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(inner_wb_o_dat[13]),
    .Z(net32),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(inner_wb_o_dat[14]),
    .Z(net33),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(inner_wb_o_dat[15]),
    .Z(net34),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(inner_wb_o_dat[1]),
    .Z(net35),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(inner_wb_o_dat[2]),
    .Z(net36),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(inner_wb_o_dat[3]),
    .Z(net37),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(inner_wb_o_dat[4]),
    .Z(net38),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(inner_wb_o_dat[5]),
    .Z(net39),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(inner_wb_adr[10]),
    .Z(net4),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(inner_wb_o_dat[6]),
    .Z(net40),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(inner_wb_o_dat[7]),
    .Z(net41),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(inner_wb_o_dat[8]),
    .Z(net42),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(inner_wb_o_dat[9]),
    .Z(net43),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(inner_wb_sel[0]),
    .Z(net44),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(inner_wb_sel[1]),
    .Z(net45),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input46 (.I(inner_wb_stb),
    .Z(net46),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input47 (.I(inner_wb_we),
    .Z(net47),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input48 (.I(iram_o_data[0]),
    .Z(net48),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input49 (.I(iram_o_data[10]),
    .Z(net49),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(inner_wb_adr[11]),
    .Z(net5),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input50 (.I(iram_o_data[11]),
    .Z(net50),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input51 (.I(iram_o_data[12]),
    .Z(net51),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(iram_o_data[13]),
    .Z(net52),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input53 (.I(iram_o_data[14]),
    .Z(net53),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input54 (.I(iram_o_data[15]),
    .Z(net54),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(iram_o_data[1]),
    .Z(net55),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(iram_o_data[2]),
    .Z(net56),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(iram_o_data[3]),
    .Z(net57),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input58 (.I(iram_o_data[4]),
    .Z(net58),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input59 (.I(iram_o_data[5]),
    .Z(net59),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(inner_wb_adr[12]),
    .Z(net6),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input60 (.I(iram_o_data[6]),
    .Z(net60),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input61 (.I(iram_o_data[7]),
    .Z(net61),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input62 (.I(iram_o_data[8]),
    .Z(net62),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input63 (.I(iram_o_data[9]),
    .Z(net63),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input64 (.I(la_data_in[0]),
    .Z(net64),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input65 (.I(la_oenb[0]),
    .Z(net65),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input66 (.I(m_io_in[0]),
    .Z(net66),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input67 (.I(m_io_in[10]),
    .Z(net67),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input68 (.I(m_io_in[11]),
    .Z(net68),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input69 (.I(m_io_in[12]),
    .Z(net69),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(inner_wb_adr[13]),
    .Z(net7),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input70 (.I(m_io_in[13]),
    .Z(net70),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input71 (.I(m_io_in[14]),
    .Z(net71),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input72 (.I(m_io_in[15]),
    .Z(net72),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input73 (.I(m_io_in[16]),
    .Z(net73),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input74 (.I(m_io_in[17]),
    .Z(net74),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input75 (.I(m_io_in[18]),
    .Z(net75),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input76 (.I(m_io_in[19]),
    .Z(net76),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input77 (.I(m_io_in[1]),
    .Z(net77),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input78 (.I(m_io_in[20]),
    .Z(net78),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input79 (.I(m_io_in[21]),
    .Z(net79),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(inner_wb_adr[14]),
    .Z(net8),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input80 (.I(m_io_in[22]),
    .Z(net80),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input81 (.I(m_io_in[23]),
    .Z(net81),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input82 (.I(m_io_in[24]),
    .Z(net82),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input83 (.I(m_io_in[25]),
    .Z(net83),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input84 (.I(m_io_in[26]),
    .Z(net84),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input85 (.I(m_io_in[27]),
    .Z(net85),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input86 (.I(m_io_in[2]),
    .Z(net86),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input87 (.I(m_io_in[30]),
    .Z(net87),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input88 (.I(m_io_in[31]),
    .Z(net88),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input89 (.I(m_io_in[32]),
    .Z(net89),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(inner_wb_adr[15]),
    .Z(net9),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input90 (.I(m_io_in[33]),
    .Z(net90),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input91 (.I(m_io_in[34]),
    .Z(net91),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input92 (.I(m_io_in[35]),
    .Z(net92),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input93 (.I(m_io_in[3]),
    .Z(net93),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input94 (.I(m_io_in[4]),
    .Z(net94),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input95 (.I(m_io_in[5]),
    .Z(net95),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input96 (.I(m_io_in[6]),
    .Z(net96),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input97 (.I(m_io_in[7]),
    .Z(net97),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input98 (.I(mgt_wb_rst_i),
    .Z(net98),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_265 (.ZN(net265),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_266 (.ZN(net266),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_267 (.ZN(net267),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_268 (.ZN(net268),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_269 (.ZN(net269),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_270 (.ZN(net270),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_271 (.ZN(net271),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_272 (.ZN(net272),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_273 (.ZN(net273),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_274 (.ZN(net274),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_275 (.ZN(net275),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_276 (.ZN(net276),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_277 (.ZN(net277),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_278 (.ZN(net278),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_279 (.ZN(net279),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_280 (.ZN(net280),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_281 (.ZN(net281),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_282 (.ZN(net282),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_283 (.ZN(net283),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_284 (.ZN(net284),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_285 (.ZN(net285),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_286 (.ZN(net286),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_287 (.ZN(net287),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_288 (.ZN(net288),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_289 (.ZN(net289),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_290 (.ZN(net290),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_291 (.ZN(net291),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_292 (.ZN(net292),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_293 (.ZN(net293),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_294 (.ZN(net294),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_295 (.ZN(net295),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_296 (.ZN(net296),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_297 (.ZN(net297),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_298 (.ZN(net298),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_299 (.ZN(net299),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_300 (.ZN(net300),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_301 (.ZN(net301),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_302 (.ZN(net302),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_303 (.ZN(net303),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_304 (.ZN(net304),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_305 (.ZN(net305),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_306 (.ZN(net306),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_307 (.ZN(net307),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_308 (.ZN(net308),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_309 (.ZN(net309),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_310 (.ZN(net310),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_311 (.ZN(net311),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_312 (.ZN(net312),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_313 (.ZN(net313),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_314 (.ZN(net314),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_315 (.ZN(net315),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_316 (.ZN(net316),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_317 (.ZN(net317),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_318 (.ZN(net318),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_319 (.ZN(net319),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_320 (.ZN(net320),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_321 (.ZN(net321),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_322 (.ZN(net322),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_323 (.ZN(net323),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_324 (.ZN(net324),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_325 (.ZN(net325),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_326 (.ZN(net326),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_327 (.ZN(net327),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_328 (.ZN(net328),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_329 (.ZN(net329),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_330 (.ZN(net330),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_331 (.ZN(net331),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_332 (.ZN(net332),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_333 (.ZN(net333),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_334 (.ZN(net334),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_335 (.ZN(net335),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_336 (.ZN(net336),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_337 (.ZN(net337),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_338 (.ZN(net338),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_339 (.ZN(net339),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_340 (.ZN(net340),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_341 (.ZN(net341),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_342 (.ZN(net342),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_343 (.ZN(net343),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_344 (.ZN(net344),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_345 (.ZN(net345),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_346 (.ZN(net346),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_347 (.ZN(net347),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_348 (.ZN(net348),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_349 (.ZN(net349),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_350 (.ZN(net350),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_351 (.ZN(net351),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_352 (.ZN(net352),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_353 (.ZN(net353),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_354 (.ZN(net354),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_355 (.ZN(net355),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_356 (.ZN(net356),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_357 (.ZN(net357),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_358 (.ZN(net358),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_359 (.ZN(net359),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_360 (.ZN(net360),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_361 (.ZN(net361),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_362 (.ZN(net362),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_363 (.ZN(net363),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_364 (.ZN(net364),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_365 (.ZN(net365),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_366 (.ZN(net366),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_367 (.ZN(net367),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_368 (.ZN(net368),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_369 (.ZN(net369),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_370 (.ZN(net370),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_371 (.ZN(net371),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_372 (.ZN(net372),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_373 (.ZN(net373),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_374 (.ZN(net374),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_375 (.ZN(net375),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_376 (.ZN(net376),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_377 (.ZN(net377),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_outer_378 (.ZN(net378),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tieh interconnect_outer_379 (.Z(net379),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tieh interconnect_outer_380 (.Z(net380),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tieh interconnect_outer_381 (.Z(net381),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tieh interconnect_outer_382 (.Z(net382),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tieh interconnect_outer_383 (.Z(net383),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tieh interconnect_outer_384 (.Z(net384),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tieh interconnect_outer_385 (.Z(net385),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tieh interconnect_outer_386 (.Z(net386),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tieh interconnect_outer_387 (.Z(net387),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap204 (.I(_1195_),
    .Z(net204),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap206 (.I(net207),
    .Z(net206),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap207 (.I(net208),
    .Z(net207),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap208 (.I(_1071_),
    .Z(net208),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 max_cap209 (.I(net210),
    .Z(net209),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 max_cap212 (.I(net213),
    .Z(net212),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 max_cap213 (.I(net214),
    .Z(net213),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap221 (.I(net222),
    .Z(net221),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap222 (.I(net223),
    .Z(net222),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap223 (.I(net224),
    .Z(net223),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap225 (.I(net226),
    .Z(net225),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap226 (.I(net227),
    .Z(net226),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap227 (.I(net228),
    .Z(net227),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap229 (.I(_0425_),
    .Z(net229),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap230 (.I(_0637_),
    .Z(net230),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap232 (.I(net233),
    .Z(net232),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap238 (.I(_1324_),
    .Z(net238),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 max_cap239 (.I(_1264_),
    .Z(net239),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 max_cap244 (.I(_0747_),
    .Z(net244),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap246 (.I(net247),
    .Z(net246),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 max_cap247 (.I(_0397_),
    .Z(net247),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap252 (.I(_1328_),
    .Z(net252),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 max_cap253 (.I(_1266_),
    .Z(net253),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap254 (.I(_1179_),
    .Z(net254),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 max_cap255 (.I(_0395_),
    .Z(net255),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap256 (.I(net257),
    .Z(net256),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap257 (.I(_1209_),
    .Z(net257),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap258 (.I(_1181_),
    .Z(net258),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 max_cap259 (.I(_0604_),
    .Z(net259),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output100 (.I(net100),
    .Z(c1_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output101 (.I(net101),
    .Z(dcache_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output102 (.I(net102),
    .Z(ic0_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output103 (.I(net103),
    .Z(ic1_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output104 (.I(net104),
    .Z(inner_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output105 (.I(net105),
    .Z(inner_disable),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output106 (.I(net106),
    .Z(inner_embed_mode),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 output107 (.I(net537),
    .Z(net391),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 output108 (.I(net392),
    .Z(net393),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output109 (.I(net109),
    .Z(inner_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output110 (.I(net110),
    .Z(inner_wb_err),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output111 (.I(net111),
    .Z(inner_wb_i_dat[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output112 (.I(net112),
    .Z(inner_wb_i_dat[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output113 (.I(net113),
    .Z(inner_wb_i_dat[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output114 (.I(net114),
    .Z(inner_wb_i_dat[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output115 (.I(net115),
    .Z(inner_wb_i_dat[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output116 (.I(net116),
    .Z(inner_wb_i_dat[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output117 (.I(net117),
    .Z(inner_wb_i_dat[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output118 (.I(net118),
    .Z(inner_wb_i_dat[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output119 (.I(net119),
    .Z(inner_wb_i_dat[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output120 (.I(net120),
    .Z(inner_wb_i_dat[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output121 (.I(net121),
    .Z(inner_wb_i_dat[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output122 (.I(net122),
    .Z(inner_wb_i_dat[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output123 (.I(net123),
    .Z(inner_wb_i_dat[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output124 (.I(net124),
    .Z(inner_wb_i_dat[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output125 (.I(net125),
    .Z(inner_wb_i_dat[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output126 (.I(net126),
    .Z(inner_wb_i_dat[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output127 (.I(net127),
    .Z(iram_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output128 (.I(net128),
    .Z(iram_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output129 (.I(net129),
    .Z(iram_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output130 (.I(net130),
    .Z(iram_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output131 (.I(net131),
    .Z(iram_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output132 (.I(net132),
    .Z(iram_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output133 (.I(net133),
    .Z(iram_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output134 (.I(net134),
    .Z(iram_i_data[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output135 (.I(net135),
    .Z(iram_i_data[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output136 (.I(net136),
    .Z(iram_i_data[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output137 (.I(net137),
    .Z(iram_i_data[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output138 (.I(net138),
    .Z(iram_i_data[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output139 (.I(net139),
    .Z(iram_i_data[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output140 (.I(net140),
    .Z(iram_i_data[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output141 (.I(net141),
    .Z(iram_i_data[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output142 (.I(net142),
    .Z(iram_i_data[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output143 (.I(net143),
    .Z(iram_i_data[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output144 (.I(net144),
    .Z(iram_i_data[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output145 (.I(net145),
    .Z(iram_i_data[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output146 (.I(net146),
    .Z(iram_i_data[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output147 (.I(net147),
    .Z(iram_i_data[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output148 (.I(net148),
    .Z(iram_i_data[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output149 (.I(net149),
    .Z(iram_i_data[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output150 (.I(net150),
    .Z(iram_we),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output151 (.I(net151),
    .Z(m_io_oeb[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output152 (.I(net152),
    .Z(m_io_oeb[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output153 (.I(net153),
    .Z(m_io_oeb[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output154 (.I(net154),
    .Z(m_io_oeb[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output155 (.I(net155),
    .Z(m_io_oeb[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output156 (.I(net156),
    .Z(m_io_oeb[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output157 (.I(net157),
    .Z(m_io_oeb[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output158 (.I(net158),
    .Z(m_io_oeb[16]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output159 (.I(net159),
    .Z(m_io_oeb[17]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output160 (.I(net160),
    .Z(m_io_oeb[18]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output161 (.I(net161),
    .Z(m_io_oeb[19]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output162 (.I(net162),
    .Z(m_io_oeb[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output163 (.I(net163),
    .Z(m_io_oeb[20]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output164 (.I(net164),
    .Z(m_io_oeb[21]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output165 (.I(net165),
    .Z(m_io_oeb[22]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output166 (.I(net166),
    .Z(m_io_oeb[23]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output167 (.I(net167),
    .Z(m_io_oeb[24]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output168 (.I(net250),
    .Z(m_io_oeb[25]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output169 (.I(net169),
    .Z(m_io_oeb[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output170 (.I(net170),
    .Z(m_io_oeb[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output171 (.I(net171),
    .Z(m_io_oeb[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output172 (.I(net172),
    .Z(m_io_oeb[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output173 (.I(net173),
    .Z(m_io_oeb[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output174 (.I(net174),
    .Z(m_io_oeb[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output175 (.I(net175),
    .Z(m_io_out[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output176 (.I(net176),
    .Z(m_io_out[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output177 (.I(net177),
    .Z(m_io_out[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output178 (.I(net178),
    .Z(m_io_out[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output179 (.I(net179),
    .Z(m_io_out[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output180 (.I(net180),
    .Z(m_io_out[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output181 (.I(net181),
    .Z(m_io_out[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output182 (.I(net182),
    .Z(m_io_out[16]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output183 (.I(net183),
    .Z(m_io_out[17]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output184 (.I(net184),
    .Z(m_io_out[18]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output185 (.I(net185),
    .Z(m_io_out[19]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output186 (.I(net186),
    .Z(m_io_out[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output187 (.I(net187),
    .Z(m_io_out[20]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output188 (.I(net188),
    .Z(m_io_out[21]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output189 (.I(net189),
    .Z(m_io_out[22]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output190 (.I(net190),
    .Z(m_io_out[23]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output191 (.I(net191),
    .Z(m_io_out[24]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output192 (.I(net192),
    .Z(m_io_out[25]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output193 (.I(net193),
    .Z(m_io_out[29]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output194 (.I(net194),
    .Z(m_io_out[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output195 (.I(net195),
    .Z(m_io_out[36]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output196 (.I(clknet_4_0_0_net196),
    .Z(m_io_out[37]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output197 (.I(net197),
    .Z(m_io_out[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output198 (.I(net198),
    .Z(m_io_out[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output199 (.I(net199),
    .Z(m_io_out[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output200 (.I(net200),
    .Z(m_io_out[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output201 (.I(net201),
    .Z(m_io_out[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output202 (.I(net202),
    .Z(m_io_out[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output203 (.I(net203),
    .Z(m_io_out[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output99 (.I(net99),
    .Z(c0_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer1 (.I(_1522_),
    .Z(net388),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer2 (.I(_1522_),
    .Z(net389),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer3 (.I(_0404_),
    .Z(net500),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire1 (.I(net495),
    .Z(net492),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire2 (.I(_1468_),
    .Z(net495),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire205 (.I(_0552_),
    .Z(net205),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 wire210 (.I(_0884_),
    .Z(net210),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 wire211 (.I(_0884_),
    .Z(net211),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 wire214 (.I(_1038_),
    .Z(net214),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire215 (.I(net525),
    .Z(net215),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire216 (.I(net519),
    .Z(net216),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire217 (.I(net522),
    .Z(net217),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire218 (.I(_0592_),
    .Z(net218),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 wire219 (.I(_0589_),
    .Z(net219),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 wire220 (.I(_1035_),
    .Z(net220),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 wire224 (.I(_0475_),
    .Z(net224),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire228 (.I(_0474_),
    .Z(net228),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 wire231 (.I(net233),
    .Z(net231),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire233 (.I(_0470_),
    .Z(net233),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire234 (.I(_1535_),
    .Z(net234),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire235 (.I(_1533_),
    .Z(net235),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire236 (.I(_1531_),
    .Z(net236),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire237 (.I(_1529_),
    .Z(net237),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 wire240 (.I(_1003_),
    .Z(net240),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire241 (.I(_1594_),
    .Z(net241),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire242 (.I(_1458_),
    .Z(net242),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 wire243 (.I(_1193_),
    .Z(net243),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire245 (.I(_0680_),
    .Z(net245),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire248 (.I(_0390_),
    .Z(net248),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire251 (.I(_1341_),
    .Z(net251),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire260 (.I(net261),
    .Z(net260),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire261 (.I(_0593_),
    .Z(net261),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire262 (.I(_0584_),
    .Z(net262),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 assign irq[0] = net265;
 assign irq[1] = net266;
 assign irq[2] = net267;
 assign la_data_out[0] = net268;
 assign la_data_out[10] = net278;
 assign la_data_out[11] = net279;
 assign la_data_out[12] = net280;
 assign la_data_out[13] = net281;
 assign la_data_out[14] = net282;
 assign la_data_out[15] = net283;
 assign la_data_out[16] = net284;
 assign la_data_out[17] = net285;
 assign la_data_out[18] = net286;
 assign la_data_out[19] = net287;
 assign la_data_out[1] = net269;
 assign la_data_out[20] = net288;
 assign la_data_out[21] = net289;
 assign la_data_out[22] = net290;
 assign la_data_out[23] = net291;
 assign la_data_out[24] = net292;
 assign la_data_out[25] = net293;
 assign la_data_out[26] = net294;
 assign la_data_out[27] = net295;
 assign la_data_out[28] = net296;
 assign la_data_out[29] = net297;
 assign la_data_out[2] = net270;
 assign la_data_out[30] = net298;
 assign la_data_out[31] = net299;
 assign la_data_out[32] = net300;
 assign la_data_out[33] = net301;
 assign la_data_out[34] = net302;
 assign la_data_out[35] = net303;
 assign la_data_out[36] = net304;
 assign la_data_out[37] = net305;
 assign la_data_out[38] = net306;
 assign la_data_out[39] = net307;
 assign la_data_out[3] = net271;
 assign la_data_out[40] = net308;
 assign la_data_out[41] = net309;
 assign la_data_out[42] = net310;
 assign la_data_out[43] = net311;
 assign la_data_out[44] = net312;
 assign la_data_out[45] = net313;
 assign la_data_out[46] = net314;
 assign la_data_out[47] = net315;
 assign la_data_out[48] = net316;
 assign la_data_out[49] = net317;
 assign la_data_out[4] = net272;
 assign la_data_out[50] = net318;
 assign la_data_out[51] = net319;
 assign la_data_out[52] = net320;
 assign la_data_out[53] = net321;
 assign la_data_out[54] = net322;
 assign la_data_out[55] = net323;
 assign la_data_out[56] = net324;
 assign la_data_out[57] = net325;
 assign la_data_out[58] = net326;
 assign la_data_out[59] = net327;
 assign la_data_out[5] = net273;
 assign la_data_out[60] = net328;
 assign la_data_out[61] = net329;
 assign la_data_out[62] = net330;
 assign la_data_out[63] = net331;
 assign la_data_out[6] = net274;
 assign la_data_out[7] = net275;
 assign la_data_out[8] = net276;
 assign la_data_out[9] = net277;
 assign m_io_oeb[26] = net379;
 assign m_io_oeb[27] = net380;
 assign m_io_oeb[28] = net334;
 assign m_io_oeb[29] = net335;
 assign m_io_oeb[30] = net381;
 assign m_io_oeb[31] = net382;
 assign m_io_oeb[32] = net383;
 assign m_io_oeb[33] = net384;
 assign m_io_oeb[34] = net385;
 assign m_io_oeb[35] = net386;
 assign m_io_oeb[36] = net336;
 assign m_io_oeb[37] = net337;
 assign m_io_oeb[8] = net332;
 assign m_io_oeb[9] = net333;
 assign m_io_out[26] = net338;
 assign m_io_out[27] = net339;
 assign m_io_out[28] = net387;
 assign m_io_out[30] = net340;
 assign m_io_out[31] = net341;
 assign m_io_out[32] = net342;
 assign m_io_out[33] = net343;
 assign m_io_out[34] = net344;
 assign m_io_out[35] = net345;
 assign mgt_wb_ack_o = net346;
 assign mgt_wb_dat_o[0] = net347;
 assign mgt_wb_dat_o[10] = net357;
 assign mgt_wb_dat_o[11] = net358;
 assign mgt_wb_dat_o[12] = net359;
 assign mgt_wb_dat_o[13] = net360;
 assign mgt_wb_dat_o[14] = net361;
 assign mgt_wb_dat_o[15] = net362;
 assign mgt_wb_dat_o[16] = net363;
 assign mgt_wb_dat_o[17] = net364;
 assign mgt_wb_dat_o[18] = net365;
 assign mgt_wb_dat_o[19] = net366;
 assign mgt_wb_dat_o[1] = net348;
 assign mgt_wb_dat_o[20] = net367;
 assign mgt_wb_dat_o[21] = net368;
 assign mgt_wb_dat_o[22] = net369;
 assign mgt_wb_dat_o[23] = net370;
 assign mgt_wb_dat_o[24] = net371;
 assign mgt_wb_dat_o[25] = net372;
 assign mgt_wb_dat_o[26] = net373;
 assign mgt_wb_dat_o[27] = net374;
 assign mgt_wb_dat_o[28] = net375;
 assign mgt_wb_dat_o[29] = net376;
 assign mgt_wb_dat_o[2] = net349;
 assign mgt_wb_dat_o[30] = net377;
 assign mgt_wb_dat_o[31] = net378;
 assign mgt_wb_dat_o[3] = net350;
 assign mgt_wb_dat_o[4] = net351;
 assign mgt_wb_dat_o[5] = net352;
 assign mgt_wb_dat_o[6] = net353;
 assign mgt_wb_dat_o[7] = net354;
 assign mgt_wb_dat_o[8] = net355;
 assign mgt_wb_dat_o[9] = net356;
endmodule
