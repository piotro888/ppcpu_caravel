magic
tech sky130A
magscale 1 2
timestamp 1672496207
<< nwell >>
rect 1066 156933 78882 157499
rect 1066 155845 78882 156411
rect 1066 154757 78882 155323
rect 1066 153669 78882 154235
rect 1066 152581 78882 153147
rect 1066 151493 78882 152059
rect 1066 150405 78882 150971
rect 1066 149317 78882 149883
rect 1066 148229 78882 148795
rect 1066 147141 78882 147707
rect 1066 146053 78882 146619
rect 1066 144965 78882 145531
rect 1066 143877 78882 144443
rect 1066 142789 78882 143355
rect 1066 141701 78882 142267
rect 1066 140613 78882 141179
rect 1066 139525 78882 140091
rect 1066 138437 78882 139003
rect 1066 137349 78882 137915
rect 1066 136261 78882 136827
rect 1066 135173 78882 135739
rect 1066 134085 78882 134651
rect 1066 132997 78882 133563
rect 1066 131909 78882 132475
rect 1066 130821 78882 131387
rect 1066 129733 78882 130299
rect 1066 128645 78882 129211
rect 1066 127557 78882 128123
rect 1066 126469 78882 127035
rect 1066 125381 78882 125947
rect 1066 124293 78882 124859
rect 1066 123205 78882 123771
rect 1066 122117 78882 122683
rect 1066 121029 78882 121595
rect 1066 119941 78882 120507
rect 1066 118853 78882 119419
rect 1066 117765 78882 118331
rect 1066 116677 78882 117243
rect 1066 115589 78882 116155
rect 1066 114501 78882 115067
rect 1066 113413 78882 113979
rect 1066 112325 78882 112891
rect 1066 111237 78882 111803
rect 1066 110149 78882 110715
rect 1066 109061 78882 109627
rect 1066 107973 78882 108539
rect 1066 106885 78882 107451
rect 1066 105797 78882 106363
rect 1066 104709 78882 105275
rect 1066 103621 78882 104187
rect 1066 102533 78882 103099
rect 1066 101445 78882 102011
rect 1066 100357 78882 100923
rect 1066 99269 78882 99835
rect 1066 98181 78882 98747
rect 1066 97093 78882 97659
rect 1066 96005 78882 96571
rect 1066 94917 78882 95483
rect 1066 93829 78882 94395
rect 1066 92741 78882 93307
rect 1066 91653 78882 92219
rect 1066 90565 78882 91131
rect 1066 89477 78882 90043
rect 1066 88389 78882 88955
rect 1066 87301 78882 87867
rect 1066 86213 78882 86779
rect 1066 85125 78882 85691
rect 1066 84037 78882 84603
rect 1066 82949 78882 83515
rect 1066 81861 78882 82427
rect 1066 80773 78882 81339
rect 1066 79685 78882 80251
rect 1066 78597 78882 79163
rect 1066 77509 78882 78075
rect 1066 76421 78882 76987
rect 1066 75333 78882 75899
rect 1066 74245 78882 74811
rect 1066 73157 78882 73723
rect 1066 72069 78882 72635
rect 1066 70981 78882 71547
rect 1066 69893 78882 70459
rect 1066 68805 78882 69371
rect 1066 67717 78882 68283
rect 1066 66629 78882 67195
rect 1066 65541 78882 66107
rect 1066 64453 78882 65019
rect 1066 63365 78882 63931
rect 1066 62277 78882 62843
rect 1066 61189 78882 61755
rect 1066 60101 78882 60667
rect 1066 59013 78882 59579
rect 1066 57925 78882 58491
rect 1066 56837 78882 57403
rect 1066 55749 78882 56315
rect 1066 54661 78882 55227
rect 1066 53573 78882 54139
rect 1066 52485 78882 53051
rect 1066 51397 78882 51963
rect 1066 50309 78882 50875
rect 1066 49221 78882 49787
rect 1066 48133 78882 48699
rect 1066 47045 78882 47611
rect 1066 45957 78882 46523
rect 1066 44869 78882 45435
rect 1066 43781 78882 44347
rect 1066 42693 78882 43259
rect 1066 41605 78882 42171
rect 1066 40517 78882 41083
rect 1066 39429 78882 39995
rect 1066 38341 78882 38907
rect 1066 37253 78882 37819
rect 1066 36165 78882 36731
rect 1066 35077 78882 35643
rect 1066 33989 78882 34555
rect 1066 32901 78882 33467
rect 1066 31813 78882 32379
rect 1066 30725 78882 31291
rect 1066 29637 78882 30203
rect 1066 28549 78882 29115
rect 1066 27461 78882 28027
rect 1066 26373 78882 26939
rect 1066 25285 78882 25851
rect 1066 24197 78882 24763
rect 1066 23109 78882 23675
rect 1066 22021 78882 22587
rect 1066 20933 78882 21499
rect 1066 19845 78882 20411
rect 1066 18757 78882 19323
rect 1066 17669 78882 18235
rect 1066 16581 78882 17147
rect 1066 15493 78882 16059
rect 1066 14405 78882 14971
rect 1066 13317 78882 13883
rect 1066 12229 78882 12795
rect 1066 11141 78882 11707
rect 1066 10053 78882 10619
rect 1066 8965 78882 9531
rect 1066 7877 78882 8443
rect 1066 6789 78882 7355
rect 1066 5701 78882 6267
rect 1066 4613 78882 5179
rect 1066 3525 78882 4091
rect 1066 2437 78882 3003
<< obsli1 >>
rect 1104 2159 78844 157777
<< obsm1 >>
rect 1104 2128 79934 157808
<< obsm2 >>
rect 4214 2139 79928 157797
<< metal3 >>
rect 79200 151648 80000 151768
rect 79200 150968 80000 151088
rect 79200 150288 80000 150408
rect 79200 149608 80000 149728
rect 79200 148928 80000 149048
rect 79200 148248 80000 148368
rect 79200 147568 80000 147688
rect 79200 146888 80000 147008
rect 79200 146208 80000 146328
rect 79200 145528 80000 145648
rect 79200 144848 80000 144968
rect 79200 144168 80000 144288
rect 79200 143488 80000 143608
rect 79200 142808 80000 142928
rect 79200 142128 80000 142248
rect 79200 141448 80000 141568
rect 79200 140768 80000 140888
rect 79200 140088 80000 140208
rect 79200 139408 80000 139528
rect 79200 138728 80000 138848
rect 79200 138048 80000 138168
rect 79200 137368 80000 137488
rect 79200 136688 80000 136808
rect 79200 136008 80000 136128
rect 79200 135328 80000 135448
rect 79200 134648 80000 134768
rect 79200 133968 80000 134088
rect 79200 133288 80000 133408
rect 79200 132608 80000 132728
rect 79200 131928 80000 132048
rect 79200 131248 80000 131368
rect 79200 130568 80000 130688
rect 79200 129888 80000 130008
rect 79200 129208 80000 129328
rect 79200 128528 80000 128648
rect 79200 127848 80000 127968
rect 79200 127168 80000 127288
rect 79200 126488 80000 126608
rect 79200 125808 80000 125928
rect 79200 125128 80000 125248
rect 79200 124448 80000 124568
rect 79200 123768 80000 123888
rect 79200 123088 80000 123208
rect 79200 122408 80000 122528
rect 79200 121728 80000 121848
rect 79200 121048 80000 121168
rect 79200 120368 80000 120488
rect 79200 119688 80000 119808
rect 79200 119008 80000 119128
rect 79200 118328 80000 118448
rect 79200 117648 80000 117768
rect 79200 116968 80000 117088
rect 79200 116288 80000 116408
rect 79200 115608 80000 115728
rect 79200 114928 80000 115048
rect 79200 114248 80000 114368
rect 79200 113568 80000 113688
rect 79200 112888 80000 113008
rect 79200 112208 80000 112328
rect 79200 111528 80000 111648
rect 79200 110848 80000 110968
rect 79200 110168 80000 110288
rect 79200 109488 80000 109608
rect 79200 108808 80000 108928
rect 79200 108128 80000 108248
rect 79200 107448 80000 107568
rect 79200 106768 80000 106888
rect 79200 106088 80000 106208
rect 79200 105408 80000 105528
rect 79200 104728 80000 104848
rect 79200 104048 80000 104168
rect 79200 103368 80000 103488
rect 79200 102688 80000 102808
rect 79200 102008 80000 102128
rect 79200 101328 80000 101448
rect 79200 100648 80000 100768
rect 79200 99968 80000 100088
rect 79200 99288 80000 99408
rect 79200 98608 80000 98728
rect 79200 97928 80000 98048
rect 79200 97248 80000 97368
rect 79200 96568 80000 96688
rect 79200 95888 80000 96008
rect 79200 95208 80000 95328
rect 79200 94528 80000 94648
rect 79200 93848 80000 93968
rect 79200 93168 80000 93288
rect 79200 92488 80000 92608
rect 79200 91808 80000 91928
rect 79200 91128 80000 91248
rect 79200 90448 80000 90568
rect 79200 89768 80000 89888
rect 79200 89088 80000 89208
rect 79200 88408 80000 88528
rect 79200 87728 80000 87848
rect 79200 87048 80000 87168
rect 79200 86368 80000 86488
rect 79200 85688 80000 85808
rect 79200 85008 80000 85128
rect 79200 84328 80000 84448
rect 79200 83648 80000 83768
rect 79200 82968 80000 83088
rect 79200 82288 80000 82408
rect 79200 81608 80000 81728
rect 79200 80928 80000 81048
rect 79200 80248 80000 80368
rect 79200 79568 80000 79688
rect 79200 78888 80000 79008
rect 79200 78208 80000 78328
rect 79200 77528 80000 77648
rect 79200 76848 80000 76968
rect 79200 76168 80000 76288
rect 79200 75488 80000 75608
rect 79200 74808 80000 74928
rect 79200 74128 80000 74248
rect 79200 73448 80000 73568
rect 79200 72768 80000 72888
rect 79200 72088 80000 72208
rect 79200 71408 80000 71528
rect 79200 70728 80000 70848
rect 79200 70048 80000 70168
rect 79200 69368 80000 69488
rect 79200 68688 80000 68808
rect 79200 68008 80000 68128
rect 79200 67328 80000 67448
rect 79200 66648 80000 66768
rect 79200 65968 80000 66088
rect 79200 65288 80000 65408
rect 79200 64608 80000 64728
rect 79200 63928 80000 64048
rect 79200 63248 80000 63368
rect 79200 62568 80000 62688
rect 79200 61888 80000 62008
rect 79200 61208 80000 61328
rect 79200 60528 80000 60648
rect 79200 59848 80000 59968
rect 79200 59168 80000 59288
rect 79200 58488 80000 58608
rect 79200 57808 80000 57928
rect 79200 57128 80000 57248
rect 79200 56448 80000 56568
rect 79200 55768 80000 55888
rect 79200 55088 80000 55208
rect 79200 54408 80000 54528
rect 79200 53728 80000 53848
rect 79200 53048 80000 53168
rect 79200 52368 80000 52488
rect 79200 51688 80000 51808
rect 79200 51008 80000 51128
rect 79200 50328 80000 50448
rect 79200 49648 80000 49768
rect 79200 48968 80000 49088
rect 79200 48288 80000 48408
rect 79200 47608 80000 47728
rect 79200 46928 80000 47048
rect 79200 46248 80000 46368
rect 79200 45568 80000 45688
rect 79200 44888 80000 45008
rect 79200 44208 80000 44328
rect 79200 43528 80000 43648
rect 79200 42848 80000 42968
rect 79200 42168 80000 42288
rect 79200 41488 80000 41608
rect 79200 40808 80000 40928
rect 79200 40128 80000 40248
rect 79200 39448 80000 39568
rect 79200 38768 80000 38888
rect 79200 38088 80000 38208
rect 79200 37408 80000 37528
rect 79200 36728 80000 36848
rect 79200 36048 80000 36168
rect 79200 35368 80000 35488
rect 79200 34688 80000 34808
rect 79200 34008 80000 34128
rect 79200 33328 80000 33448
rect 79200 32648 80000 32768
rect 79200 31968 80000 32088
rect 79200 31288 80000 31408
rect 79200 30608 80000 30728
rect 79200 29928 80000 30048
rect 79200 29248 80000 29368
rect 79200 28568 80000 28688
rect 79200 27888 80000 28008
rect 79200 27208 80000 27328
rect 79200 26528 80000 26648
rect 79200 25848 80000 25968
rect 79200 25168 80000 25288
rect 79200 24488 80000 24608
rect 79200 23808 80000 23928
rect 79200 23128 80000 23248
rect 79200 22448 80000 22568
rect 79200 21768 80000 21888
rect 79200 21088 80000 21208
rect 79200 20408 80000 20528
rect 79200 19728 80000 19848
rect 79200 19048 80000 19168
rect 79200 18368 80000 18488
rect 79200 17688 80000 17808
rect 79200 17008 80000 17128
rect 79200 16328 80000 16448
rect 79200 15648 80000 15768
rect 79200 14968 80000 15088
rect 79200 14288 80000 14408
rect 79200 13608 80000 13728
rect 79200 12928 80000 13048
rect 79200 12248 80000 12368
rect 79200 11568 80000 11688
rect 79200 10888 80000 11008
rect 79200 10208 80000 10328
rect 79200 9528 80000 9648
rect 79200 8848 80000 8968
rect 79200 8168 80000 8288
<< obsm3 >>
rect 4210 151848 79200 157793
rect 4210 151568 79120 151848
rect 4210 151168 79200 151568
rect 4210 150888 79120 151168
rect 4210 150488 79200 150888
rect 4210 150208 79120 150488
rect 4210 149808 79200 150208
rect 4210 149528 79120 149808
rect 4210 149128 79200 149528
rect 4210 148848 79120 149128
rect 4210 148448 79200 148848
rect 4210 148168 79120 148448
rect 4210 147768 79200 148168
rect 4210 147488 79120 147768
rect 4210 147088 79200 147488
rect 4210 146808 79120 147088
rect 4210 146408 79200 146808
rect 4210 146128 79120 146408
rect 4210 145728 79200 146128
rect 4210 145448 79120 145728
rect 4210 145048 79200 145448
rect 4210 144768 79120 145048
rect 4210 144368 79200 144768
rect 4210 144088 79120 144368
rect 4210 143688 79200 144088
rect 4210 143408 79120 143688
rect 4210 143008 79200 143408
rect 4210 142728 79120 143008
rect 4210 142328 79200 142728
rect 4210 142048 79120 142328
rect 4210 141648 79200 142048
rect 4210 141368 79120 141648
rect 4210 140968 79200 141368
rect 4210 140688 79120 140968
rect 4210 140288 79200 140688
rect 4210 140008 79120 140288
rect 4210 139608 79200 140008
rect 4210 139328 79120 139608
rect 4210 138928 79200 139328
rect 4210 138648 79120 138928
rect 4210 138248 79200 138648
rect 4210 137968 79120 138248
rect 4210 137568 79200 137968
rect 4210 137288 79120 137568
rect 4210 136888 79200 137288
rect 4210 136608 79120 136888
rect 4210 136208 79200 136608
rect 4210 135928 79120 136208
rect 4210 135528 79200 135928
rect 4210 135248 79120 135528
rect 4210 134848 79200 135248
rect 4210 134568 79120 134848
rect 4210 134168 79200 134568
rect 4210 133888 79120 134168
rect 4210 133488 79200 133888
rect 4210 133208 79120 133488
rect 4210 132808 79200 133208
rect 4210 132528 79120 132808
rect 4210 132128 79200 132528
rect 4210 131848 79120 132128
rect 4210 131448 79200 131848
rect 4210 131168 79120 131448
rect 4210 130768 79200 131168
rect 4210 130488 79120 130768
rect 4210 130088 79200 130488
rect 4210 129808 79120 130088
rect 4210 129408 79200 129808
rect 4210 129128 79120 129408
rect 4210 128728 79200 129128
rect 4210 128448 79120 128728
rect 4210 128048 79200 128448
rect 4210 127768 79120 128048
rect 4210 127368 79200 127768
rect 4210 127088 79120 127368
rect 4210 126688 79200 127088
rect 4210 126408 79120 126688
rect 4210 126008 79200 126408
rect 4210 125728 79120 126008
rect 4210 125328 79200 125728
rect 4210 125048 79120 125328
rect 4210 124648 79200 125048
rect 4210 124368 79120 124648
rect 4210 123968 79200 124368
rect 4210 123688 79120 123968
rect 4210 123288 79200 123688
rect 4210 123008 79120 123288
rect 4210 122608 79200 123008
rect 4210 122328 79120 122608
rect 4210 121928 79200 122328
rect 4210 121648 79120 121928
rect 4210 121248 79200 121648
rect 4210 120968 79120 121248
rect 4210 120568 79200 120968
rect 4210 120288 79120 120568
rect 4210 119888 79200 120288
rect 4210 119608 79120 119888
rect 4210 119208 79200 119608
rect 4210 118928 79120 119208
rect 4210 118528 79200 118928
rect 4210 118248 79120 118528
rect 4210 117848 79200 118248
rect 4210 117568 79120 117848
rect 4210 117168 79200 117568
rect 4210 116888 79120 117168
rect 4210 116488 79200 116888
rect 4210 116208 79120 116488
rect 4210 115808 79200 116208
rect 4210 115528 79120 115808
rect 4210 115128 79200 115528
rect 4210 114848 79120 115128
rect 4210 114448 79200 114848
rect 4210 114168 79120 114448
rect 4210 113768 79200 114168
rect 4210 113488 79120 113768
rect 4210 113088 79200 113488
rect 4210 112808 79120 113088
rect 4210 112408 79200 112808
rect 4210 112128 79120 112408
rect 4210 111728 79200 112128
rect 4210 111448 79120 111728
rect 4210 111048 79200 111448
rect 4210 110768 79120 111048
rect 4210 110368 79200 110768
rect 4210 110088 79120 110368
rect 4210 109688 79200 110088
rect 4210 109408 79120 109688
rect 4210 109008 79200 109408
rect 4210 108728 79120 109008
rect 4210 108328 79200 108728
rect 4210 108048 79120 108328
rect 4210 107648 79200 108048
rect 4210 107368 79120 107648
rect 4210 106968 79200 107368
rect 4210 106688 79120 106968
rect 4210 106288 79200 106688
rect 4210 106008 79120 106288
rect 4210 105608 79200 106008
rect 4210 105328 79120 105608
rect 4210 104928 79200 105328
rect 4210 104648 79120 104928
rect 4210 104248 79200 104648
rect 4210 103968 79120 104248
rect 4210 103568 79200 103968
rect 4210 103288 79120 103568
rect 4210 102888 79200 103288
rect 4210 102608 79120 102888
rect 4210 102208 79200 102608
rect 4210 101928 79120 102208
rect 4210 101528 79200 101928
rect 4210 101248 79120 101528
rect 4210 100848 79200 101248
rect 4210 100568 79120 100848
rect 4210 100168 79200 100568
rect 4210 99888 79120 100168
rect 4210 99488 79200 99888
rect 4210 99208 79120 99488
rect 4210 98808 79200 99208
rect 4210 98528 79120 98808
rect 4210 98128 79200 98528
rect 4210 97848 79120 98128
rect 4210 97448 79200 97848
rect 4210 97168 79120 97448
rect 4210 96768 79200 97168
rect 4210 96488 79120 96768
rect 4210 96088 79200 96488
rect 4210 95808 79120 96088
rect 4210 95408 79200 95808
rect 4210 95128 79120 95408
rect 4210 94728 79200 95128
rect 4210 94448 79120 94728
rect 4210 94048 79200 94448
rect 4210 93768 79120 94048
rect 4210 93368 79200 93768
rect 4210 93088 79120 93368
rect 4210 92688 79200 93088
rect 4210 92408 79120 92688
rect 4210 92008 79200 92408
rect 4210 91728 79120 92008
rect 4210 91328 79200 91728
rect 4210 91048 79120 91328
rect 4210 90648 79200 91048
rect 4210 90368 79120 90648
rect 4210 89968 79200 90368
rect 4210 89688 79120 89968
rect 4210 89288 79200 89688
rect 4210 89008 79120 89288
rect 4210 88608 79200 89008
rect 4210 88328 79120 88608
rect 4210 87928 79200 88328
rect 4210 87648 79120 87928
rect 4210 87248 79200 87648
rect 4210 86968 79120 87248
rect 4210 86568 79200 86968
rect 4210 86288 79120 86568
rect 4210 85888 79200 86288
rect 4210 85608 79120 85888
rect 4210 85208 79200 85608
rect 4210 84928 79120 85208
rect 4210 84528 79200 84928
rect 4210 84248 79120 84528
rect 4210 83848 79200 84248
rect 4210 83568 79120 83848
rect 4210 83168 79200 83568
rect 4210 82888 79120 83168
rect 4210 82488 79200 82888
rect 4210 82208 79120 82488
rect 4210 81808 79200 82208
rect 4210 81528 79120 81808
rect 4210 81128 79200 81528
rect 4210 80848 79120 81128
rect 4210 80448 79200 80848
rect 4210 80168 79120 80448
rect 4210 79768 79200 80168
rect 4210 79488 79120 79768
rect 4210 79088 79200 79488
rect 4210 78808 79120 79088
rect 4210 78408 79200 78808
rect 4210 78128 79120 78408
rect 4210 77728 79200 78128
rect 4210 77448 79120 77728
rect 4210 77048 79200 77448
rect 4210 76768 79120 77048
rect 4210 76368 79200 76768
rect 4210 76088 79120 76368
rect 4210 75688 79200 76088
rect 4210 75408 79120 75688
rect 4210 75008 79200 75408
rect 4210 74728 79120 75008
rect 4210 74328 79200 74728
rect 4210 74048 79120 74328
rect 4210 73648 79200 74048
rect 4210 73368 79120 73648
rect 4210 72968 79200 73368
rect 4210 72688 79120 72968
rect 4210 72288 79200 72688
rect 4210 72008 79120 72288
rect 4210 71608 79200 72008
rect 4210 71328 79120 71608
rect 4210 70928 79200 71328
rect 4210 70648 79120 70928
rect 4210 70248 79200 70648
rect 4210 69968 79120 70248
rect 4210 69568 79200 69968
rect 4210 69288 79120 69568
rect 4210 68888 79200 69288
rect 4210 68608 79120 68888
rect 4210 68208 79200 68608
rect 4210 67928 79120 68208
rect 4210 67528 79200 67928
rect 4210 67248 79120 67528
rect 4210 66848 79200 67248
rect 4210 66568 79120 66848
rect 4210 66168 79200 66568
rect 4210 65888 79120 66168
rect 4210 65488 79200 65888
rect 4210 65208 79120 65488
rect 4210 64808 79200 65208
rect 4210 64528 79120 64808
rect 4210 64128 79200 64528
rect 4210 63848 79120 64128
rect 4210 63448 79200 63848
rect 4210 63168 79120 63448
rect 4210 62768 79200 63168
rect 4210 62488 79120 62768
rect 4210 62088 79200 62488
rect 4210 61808 79120 62088
rect 4210 61408 79200 61808
rect 4210 61128 79120 61408
rect 4210 60728 79200 61128
rect 4210 60448 79120 60728
rect 4210 60048 79200 60448
rect 4210 59768 79120 60048
rect 4210 59368 79200 59768
rect 4210 59088 79120 59368
rect 4210 58688 79200 59088
rect 4210 58408 79120 58688
rect 4210 58008 79200 58408
rect 4210 57728 79120 58008
rect 4210 57328 79200 57728
rect 4210 57048 79120 57328
rect 4210 56648 79200 57048
rect 4210 56368 79120 56648
rect 4210 55968 79200 56368
rect 4210 55688 79120 55968
rect 4210 55288 79200 55688
rect 4210 55008 79120 55288
rect 4210 54608 79200 55008
rect 4210 54328 79120 54608
rect 4210 53928 79200 54328
rect 4210 53648 79120 53928
rect 4210 53248 79200 53648
rect 4210 52968 79120 53248
rect 4210 52568 79200 52968
rect 4210 52288 79120 52568
rect 4210 51888 79200 52288
rect 4210 51608 79120 51888
rect 4210 51208 79200 51608
rect 4210 50928 79120 51208
rect 4210 50528 79200 50928
rect 4210 50248 79120 50528
rect 4210 49848 79200 50248
rect 4210 49568 79120 49848
rect 4210 49168 79200 49568
rect 4210 48888 79120 49168
rect 4210 48488 79200 48888
rect 4210 48208 79120 48488
rect 4210 47808 79200 48208
rect 4210 47528 79120 47808
rect 4210 47128 79200 47528
rect 4210 46848 79120 47128
rect 4210 46448 79200 46848
rect 4210 46168 79120 46448
rect 4210 45768 79200 46168
rect 4210 45488 79120 45768
rect 4210 45088 79200 45488
rect 4210 44808 79120 45088
rect 4210 44408 79200 44808
rect 4210 44128 79120 44408
rect 4210 43728 79200 44128
rect 4210 43448 79120 43728
rect 4210 43048 79200 43448
rect 4210 42768 79120 43048
rect 4210 42368 79200 42768
rect 4210 42088 79120 42368
rect 4210 41688 79200 42088
rect 4210 41408 79120 41688
rect 4210 41008 79200 41408
rect 4210 40728 79120 41008
rect 4210 40328 79200 40728
rect 4210 40048 79120 40328
rect 4210 39648 79200 40048
rect 4210 39368 79120 39648
rect 4210 38968 79200 39368
rect 4210 38688 79120 38968
rect 4210 38288 79200 38688
rect 4210 38008 79120 38288
rect 4210 37608 79200 38008
rect 4210 37328 79120 37608
rect 4210 36928 79200 37328
rect 4210 36648 79120 36928
rect 4210 36248 79200 36648
rect 4210 35968 79120 36248
rect 4210 35568 79200 35968
rect 4210 35288 79120 35568
rect 4210 34888 79200 35288
rect 4210 34608 79120 34888
rect 4210 34208 79200 34608
rect 4210 33928 79120 34208
rect 4210 33528 79200 33928
rect 4210 33248 79120 33528
rect 4210 32848 79200 33248
rect 4210 32568 79120 32848
rect 4210 32168 79200 32568
rect 4210 31888 79120 32168
rect 4210 31488 79200 31888
rect 4210 31208 79120 31488
rect 4210 30808 79200 31208
rect 4210 30528 79120 30808
rect 4210 30128 79200 30528
rect 4210 29848 79120 30128
rect 4210 29448 79200 29848
rect 4210 29168 79120 29448
rect 4210 28768 79200 29168
rect 4210 28488 79120 28768
rect 4210 28088 79200 28488
rect 4210 27808 79120 28088
rect 4210 27408 79200 27808
rect 4210 27128 79120 27408
rect 4210 26728 79200 27128
rect 4210 26448 79120 26728
rect 4210 26048 79200 26448
rect 4210 25768 79120 26048
rect 4210 25368 79200 25768
rect 4210 25088 79120 25368
rect 4210 24688 79200 25088
rect 4210 24408 79120 24688
rect 4210 24008 79200 24408
rect 4210 23728 79120 24008
rect 4210 23328 79200 23728
rect 4210 23048 79120 23328
rect 4210 22648 79200 23048
rect 4210 22368 79120 22648
rect 4210 21968 79200 22368
rect 4210 21688 79120 21968
rect 4210 21288 79200 21688
rect 4210 21008 79120 21288
rect 4210 20608 79200 21008
rect 4210 20328 79120 20608
rect 4210 19928 79200 20328
rect 4210 19648 79120 19928
rect 4210 19248 79200 19648
rect 4210 18968 79120 19248
rect 4210 18568 79200 18968
rect 4210 18288 79120 18568
rect 4210 17888 79200 18288
rect 4210 17608 79120 17888
rect 4210 17208 79200 17608
rect 4210 16928 79120 17208
rect 4210 16528 79200 16928
rect 4210 16248 79120 16528
rect 4210 15848 79200 16248
rect 4210 15568 79120 15848
rect 4210 15168 79200 15568
rect 4210 14888 79120 15168
rect 4210 14488 79200 14888
rect 4210 14208 79120 14488
rect 4210 13808 79200 14208
rect 4210 13528 79120 13808
rect 4210 13128 79200 13528
rect 4210 12848 79120 13128
rect 4210 12448 79200 12848
rect 4210 12168 79120 12448
rect 4210 11768 79200 12168
rect 4210 11488 79120 11768
rect 4210 11088 79200 11488
rect 4210 10808 79120 11088
rect 4210 10408 79200 10808
rect 4210 10128 79120 10408
rect 4210 9728 79200 10128
rect 4210 9448 79120 9728
rect 4210 9048 79200 9448
rect 4210 8768 79120 9048
rect 4210 8368 79200 8768
rect 4210 8088 79120 8368
rect 4210 2143 79200 8088
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
<< obsm4 >>
rect 34467 9555 34848 153645
rect 35328 9555 50208 153645
rect 50688 9555 65568 153645
rect 66048 9555 77221 153645
<< labels >>
rlabel metal3 s 79200 20408 80000 20528 6 dbg_pc[0]
port 1 nsew signal output
rlabel metal3 s 79200 100648 80000 100768 6 dbg_pc[10]
port 2 nsew signal output
rlabel metal3 s 79200 107448 80000 107568 6 dbg_pc[11]
port 3 nsew signal output
rlabel metal3 s 79200 114248 80000 114368 6 dbg_pc[12]
port 4 nsew signal output
rlabel metal3 s 79200 121048 80000 121168 6 dbg_pc[13]
port 5 nsew signal output
rlabel metal3 s 79200 127848 80000 127968 6 dbg_pc[14]
port 6 nsew signal output
rlabel metal3 s 79200 134648 80000 134768 6 dbg_pc[15]
port 7 nsew signal output
rlabel metal3 s 79200 29248 80000 29368 6 dbg_pc[1]
port 8 nsew signal output
rlabel metal3 s 79200 38088 80000 38208 6 dbg_pc[2]
port 9 nsew signal output
rlabel metal3 s 79200 46248 80000 46368 6 dbg_pc[3]
port 10 nsew signal output
rlabel metal3 s 79200 54408 80000 54528 6 dbg_pc[4]
port 11 nsew signal output
rlabel metal3 s 79200 62568 80000 62688 6 dbg_pc[5]
port 12 nsew signal output
rlabel metal3 s 79200 70728 80000 70848 6 dbg_pc[6]
port 13 nsew signal output
rlabel metal3 s 79200 78888 80000 79008 6 dbg_pc[7]
port 14 nsew signal output
rlabel metal3 s 79200 87048 80000 87168 6 dbg_pc[8]
port 15 nsew signal output
rlabel metal3 s 79200 93848 80000 93968 6 dbg_pc[9]
port 16 nsew signal output
rlabel metal3 s 79200 21088 80000 21208 6 dbg_r0[0]
port 17 nsew signal output
rlabel metal3 s 79200 101328 80000 101448 6 dbg_r0[10]
port 18 nsew signal output
rlabel metal3 s 79200 108128 80000 108248 6 dbg_r0[11]
port 19 nsew signal output
rlabel metal3 s 79200 114928 80000 115048 6 dbg_r0[12]
port 20 nsew signal output
rlabel metal3 s 79200 121728 80000 121848 6 dbg_r0[13]
port 21 nsew signal output
rlabel metal3 s 79200 128528 80000 128648 6 dbg_r0[14]
port 22 nsew signal output
rlabel metal3 s 79200 135328 80000 135448 6 dbg_r0[15]
port 23 nsew signal output
rlabel metal3 s 79200 29928 80000 30048 6 dbg_r0[1]
port 24 nsew signal output
rlabel metal3 s 79200 38768 80000 38888 6 dbg_r0[2]
port 25 nsew signal output
rlabel metal3 s 79200 46928 80000 47048 6 dbg_r0[3]
port 26 nsew signal output
rlabel metal3 s 79200 55088 80000 55208 6 dbg_r0[4]
port 27 nsew signal output
rlabel metal3 s 79200 63248 80000 63368 6 dbg_r0[5]
port 28 nsew signal output
rlabel metal3 s 79200 71408 80000 71528 6 dbg_r0[6]
port 29 nsew signal output
rlabel metal3 s 79200 79568 80000 79688 6 dbg_r0[7]
port 30 nsew signal output
rlabel metal3 s 79200 87728 80000 87848 6 dbg_r0[8]
port 31 nsew signal output
rlabel metal3 s 79200 94528 80000 94648 6 dbg_r0[9]
port 32 nsew signal output
rlabel metal3 s 79200 8168 80000 8288 6 i_clk
port 33 nsew signal input
rlabel metal3 s 79200 21768 80000 21888 6 i_core_int_sreg[0]
port 34 nsew signal input
rlabel metal3 s 79200 102008 80000 102128 6 i_core_int_sreg[10]
port 35 nsew signal input
rlabel metal3 s 79200 108808 80000 108928 6 i_core_int_sreg[11]
port 36 nsew signal input
rlabel metal3 s 79200 115608 80000 115728 6 i_core_int_sreg[12]
port 37 nsew signal input
rlabel metal3 s 79200 122408 80000 122528 6 i_core_int_sreg[13]
port 38 nsew signal input
rlabel metal3 s 79200 129208 80000 129328 6 i_core_int_sreg[14]
port 39 nsew signal input
rlabel metal3 s 79200 136008 80000 136128 6 i_core_int_sreg[15]
port 40 nsew signal input
rlabel metal3 s 79200 30608 80000 30728 6 i_core_int_sreg[1]
port 41 nsew signal input
rlabel metal3 s 79200 39448 80000 39568 6 i_core_int_sreg[2]
port 42 nsew signal input
rlabel metal3 s 79200 47608 80000 47728 6 i_core_int_sreg[3]
port 43 nsew signal input
rlabel metal3 s 79200 55768 80000 55888 6 i_core_int_sreg[4]
port 44 nsew signal input
rlabel metal3 s 79200 63928 80000 64048 6 i_core_int_sreg[5]
port 45 nsew signal input
rlabel metal3 s 79200 72088 80000 72208 6 i_core_int_sreg[6]
port 46 nsew signal input
rlabel metal3 s 79200 80248 80000 80368 6 i_core_int_sreg[7]
port 47 nsew signal input
rlabel metal3 s 79200 88408 80000 88528 6 i_core_int_sreg[8]
port 48 nsew signal input
rlabel metal3 s 79200 95208 80000 95328 6 i_core_int_sreg[9]
port 49 nsew signal input
rlabel metal3 s 79200 8848 80000 8968 6 i_disable
port 50 nsew signal input
rlabel metal3 s 79200 9528 80000 9648 6 i_irq
port 51 nsew signal input
rlabel metal3 s 79200 10208 80000 10328 6 i_mc_core_int
port 52 nsew signal input
rlabel metal3 s 79200 10888 80000 11008 6 i_mem_ack
port 53 nsew signal input
rlabel metal3 s 79200 22448 80000 22568 6 i_mem_data[0]
port 54 nsew signal input
rlabel metal3 s 79200 102688 80000 102808 6 i_mem_data[10]
port 55 nsew signal input
rlabel metal3 s 79200 109488 80000 109608 6 i_mem_data[11]
port 56 nsew signal input
rlabel metal3 s 79200 116288 80000 116408 6 i_mem_data[12]
port 57 nsew signal input
rlabel metal3 s 79200 123088 80000 123208 6 i_mem_data[13]
port 58 nsew signal input
rlabel metal3 s 79200 129888 80000 130008 6 i_mem_data[14]
port 59 nsew signal input
rlabel metal3 s 79200 136688 80000 136808 6 i_mem_data[15]
port 60 nsew signal input
rlabel metal3 s 79200 31288 80000 31408 6 i_mem_data[1]
port 61 nsew signal input
rlabel metal3 s 79200 40128 80000 40248 6 i_mem_data[2]
port 62 nsew signal input
rlabel metal3 s 79200 48288 80000 48408 6 i_mem_data[3]
port 63 nsew signal input
rlabel metal3 s 79200 56448 80000 56568 6 i_mem_data[4]
port 64 nsew signal input
rlabel metal3 s 79200 64608 80000 64728 6 i_mem_data[5]
port 65 nsew signal input
rlabel metal3 s 79200 72768 80000 72888 6 i_mem_data[6]
port 66 nsew signal input
rlabel metal3 s 79200 80928 80000 81048 6 i_mem_data[7]
port 67 nsew signal input
rlabel metal3 s 79200 89088 80000 89208 6 i_mem_data[8]
port 68 nsew signal input
rlabel metal3 s 79200 95888 80000 96008 6 i_mem_data[9]
port 69 nsew signal input
rlabel metal3 s 79200 11568 80000 11688 6 i_mem_exception
port 70 nsew signal input
rlabel metal3 s 79200 23128 80000 23248 6 i_req_data[0]
port 71 nsew signal input
rlabel metal3 s 79200 103368 80000 103488 6 i_req_data[10]
port 72 nsew signal input
rlabel metal3 s 79200 110168 80000 110288 6 i_req_data[11]
port 73 nsew signal input
rlabel metal3 s 79200 116968 80000 117088 6 i_req_data[12]
port 74 nsew signal input
rlabel metal3 s 79200 123768 80000 123888 6 i_req_data[13]
port 75 nsew signal input
rlabel metal3 s 79200 130568 80000 130688 6 i_req_data[14]
port 76 nsew signal input
rlabel metal3 s 79200 137368 80000 137488 6 i_req_data[15]
port 77 nsew signal input
rlabel metal3 s 79200 141448 80000 141568 6 i_req_data[16]
port 78 nsew signal input
rlabel metal3 s 79200 142128 80000 142248 6 i_req_data[17]
port 79 nsew signal input
rlabel metal3 s 79200 142808 80000 142928 6 i_req_data[18]
port 80 nsew signal input
rlabel metal3 s 79200 143488 80000 143608 6 i_req_data[19]
port 81 nsew signal input
rlabel metal3 s 79200 31968 80000 32088 6 i_req_data[1]
port 82 nsew signal input
rlabel metal3 s 79200 144168 80000 144288 6 i_req_data[20]
port 83 nsew signal input
rlabel metal3 s 79200 144848 80000 144968 6 i_req_data[21]
port 84 nsew signal input
rlabel metal3 s 79200 145528 80000 145648 6 i_req_data[22]
port 85 nsew signal input
rlabel metal3 s 79200 146208 80000 146328 6 i_req_data[23]
port 86 nsew signal input
rlabel metal3 s 79200 146888 80000 147008 6 i_req_data[24]
port 87 nsew signal input
rlabel metal3 s 79200 147568 80000 147688 6 i_req_data[25]
port 88 nsew signal input
rlabel metal3 s 79200 148248 80000 148368 6 i_req_data[26]
port 89 nsew signal input
rlabel metal3 s 79200 148928 80000 149048 6 i_req_data[27]
port 90 nsew signal input
rlabel metal3 s 79200 149608 80000 149728 6 i_req_data[28]
port 91 nsew signal input
rlabel metal3 s 79200 150288 80000 150408 6 i_req_data[29]
port 92 nsew signal input
rlabel metal3 s 79200 40808 80000 40928 6 i_req_data[2]
port 93 nsew signal input
rlabel metal3 s 79200 150968 80000 151088 6 i_req_data[30]
port 94 nsew signal input
rlabel metal3 s 79200 151648 80000 151768 6 i_req_data[31]
port 95 nsew signal input
rlabel metal3 s 79200 48968 80000 49088 6 i_req_data[3]
port 96 nsew signal input
rlabel metal3 s 79200 57128 80000 57248 6 i_req_data[4]
port 97 nsew signal input
rlabel metal3 s 79200 65288 80000 65408 6 i_req_data[5]
port 98 nsew signal input
rlabel metal3 s 79200 73448 80000 73568 6 i_req_data[6]
port 99 nsew signal input
rlabel metal3 s 79200 81608 80000 81728 6 i_req_data[7]
port 100 nsew signal input
rlabel metal3 s 79200 89768 80000 89888 6 i_req_data[8]
port 101 nsew signal input
rlabel metal3 s 79200 96568 80000 96688 6 i_req_data[9]
port 102 nsew signal input
rlabel metal3 s 79200 12248 80000 12368 6 i_req_data_valid
port 103 nsew signal input
rlabel metal3 s 79200 12928 80000 13048 6 i_rst
port 104 nsew signal input
rlabel metal3 s 79200 13608 80000 13728 6 o_c_data_page
port 105 nsew signal output
rlabel metal3 s 79200 14288 80000 14408 6 o_c_instr_long
port 106 nsew signal output
rlabel metal3 s 79200 14968 80000 15088 6 o_c_instr_page
port 107 nsew signal output
rlabel metal3 s 79200 15648 80000 15768 6 o_icache_flush
port 108 nsew signal output
rlabel metal3 s 79200 23808 80000 23928 6 o_instr_long_addr[0]
port 109 nsew signal output
rlabel metal3 s 79200 32648 80000 32768 6 o_instr_long_addr[1]
port 110 nsew signal output
rlabel metal3 s 79200 41488 80000 41608 6 o_instr_long_addr[2]
port 111 nsew signal output
rlabel metal3 s 79200 49648 80000 49768 6 o_instr_long_addr[3]
port 112 nsew signal output
rlabel metal3 s 79200 57808 80000 57928 6 o_instr_long_addr[4]
port 113 nsew signal output
rlabel metal3 s 79200 65968 80000 66088 6 o_instr_long_addr[5]
port 114 nsew signal output
rlabel metal3 s 79200 74128 80000 74248 6 o_instr_long_addr[6]
port 115 nsew signal output
rlabel metal3 s 79200 82288 80000 82408 6 o_instr_long_addr[7]
port 116 nsew signal output
rlabel metal3 s 79200 24488 80000 24608 6 o_mem_addr[0]
port 117 nsew signal output
rlabel metal3 s 79200 104048 80000 104168 6 o_mem_addr[10]
port 118 nsew signal output
rlabel metal3 s 79200 110848 80000 110968 6 o_mem_addr[11]
port 119 nsew signal output
rlabel metal3 s 79200 117648 80000 117768 6 o_mem_addr[12]
port 120 nsew signal output
rlabel metal3 s 79200 124448 80000 124568 6 o_mem_addr[13]
port 121 nsew signal output
rlabel metal3 s 79200 131248 80000 131368 6 o_mem_addr[14]
port 122 nsew signal output
rlabel metal3 s 79200 138048 80000 138168 6 o_mem_addr[15]
port 123 nsew signal output
rlabel metal3 s 79200 33328 80000 33448 6 o_mem_addr[1]
port 124 nsew signal output
rlabel metal3 s 79200 42168 80000 42288 6 o_mem_addr[2]
port 125 nsew signal output
rlabel metal3 s 79200 50328 80000 50448 6 o_mem_addr[3]
port 126 nsew signal output
rlabel metal3 s 79200 58488 80000 58608 6 o_mem_addr[4]
port 127 nsew signal output
rlabel metal3 s 79200 66648 80000 66768 6 o_mem_addr[5]
port 128 nsew signal output
rlabel metal3 s 79200 74808 80000 74928 6 o_mem_addr[6]
port 129 nsew signal output
rlabel metal3 s 79200 82968 80000 83088 6 o_mem_addr[7]
port 130 nsew signal output
rlabel metal3 s 79200 90448 80000 90568 6 o_mem_addr[8]
port 131 nsew signal output
rlabel metal3 s 79200 97248 80000 97368 6 o_mem_addr[9]
port 132 nsew signal output
rlabel metal3 s 79200 25168 80000 25288 6 o_mem_addr_high[0]
port 133 nsew signal output
rlabel metal3 s 79200 34008 80000 34128 6 o_mem_addr_high[1]
port 134 nsew signal output
rlabel metal3 s 79200 42848 80000 42968 6 o_mem_addr_high[2]
port 135 nsew signal output
rlabel metal3 s 79200 51008 80000 51128 6 o_mem_addr_high[3]
port 136 nsew signal output
rlabel metal3 s 79200 59168 80000 59288 6 o_mem_addr_high[4]
port 137 nsew signal output
rlabel metal3 s 79200 67328 80000 67448 6 o_mem_addr_high[5]
port 138 nsew signal output
rlabel metal3 s 79200 75488 80000 75608 6 o_mem_addr_high[6]
port 139 nsew signal output
rlabel metal3 s 79200 83648 80000 83768 6 o_mem_addr_high[7]
port 140 nsew signal output
rlabel metal3 s 79200 25848 80000 25968 6 o_mem_data[0]
port 141 nsew signal output
rlabel metal3 s 79200 104728 80000 104848 6 o_mem_data[10]
port 142 nsew signal output
rlabel metal3 s 79200 111528 80000 111648 6 o_mem_data[11]
port 143 nsew signal output
rlabel metal3 s 79200 118328 80000 118448 6 o_mem_data[12]
port 144 nsew signal output
rlabel metal3 s 79200 125128 80000 125248 6 o_mem_data[13]
port 145 nsew signal output
rlabel metal3 s 79200 131928 80000 132048 6 o_mem_data[14]
port 146 nsew signal output
rlabel metal3 s 79200 138728 80000 138848 6 o_mem_data[15]
port 147 nsew signal output
rlabel metal3 s 79200 34688 80000 34808 6 o_mem_data[1]
port 148 nsew signal output
rlabel metal3 s 79200 43528 80000 43648 6 o_mem_data[2]
port 149 nsew signal output
rlabel metal3 s 79200 51688 80000 51808 6 o_mem_data[3]
port 150 nsew signal output
rlabel metal3 s 79200 59848 80000 59968 6 o_mem_data[4]
port 151 nsew signal output
rlabel metal3 s 79200 68008 80000 68128 6 o_mem_data[5]
port 152 nsew signal output
rlabel metal3 s 79200 76168 80000 76288 6 o_mem_data[6]
port 153 nsew signal output
rlabel metal3 s 79200 84328 80000 84448 6 o_mem_data[7]
port 154 nsew signal output
rlabel metal3 s 79200 91128 80000 91248 6 o_mem_data[8]
port 155 nsew signal output
rlabel metal3 s 79200 97928 80000 98048 6 o_mem_data[9]
port 156 nsew signal output
rlabel metal3 s 79200 16328 80000 16448 6 o_mem_long
port 157 nsew signal output
rlabel metal3 s 79200 17008 80000 17128 6 o_mem_req
port 158 nsew signal output
rlabel metal3 s 79200 26528 80000 26648 6 o_mem_sel[0]
port 159 nsew signal output
rlabel metal3 s 79200 35368 80000 35488 6 o_mem_sel[1]
port 160 nsew signal output
rlabel metal3 s 79200 17688 80000 17808 6 o_mem_we
port 161 nsew signal output
rlabel metal3 s 79200 18368 80000 18488 6 o_req_active
port 162 nsew signal output
rlabel metal3 s 79200 27208 80000 27328 6 o_req_addr[0]
port 163 nsew signal output
rlabel metal3 s 79200 105408 80000 105528 6 o_req_addr[10]
port 164 nsew signal output
rlabel metal3 s 79200 112208 80000 112328 6 o_req_addr[11]
port 165 nsew signal output
rlabel metal3 s 79200 119008 80000 119128 6 o_req_addr[12]
port 166 nsew signal output
rlabel metal3 s 79200 125808 80000 125928 6 o_req_addr[13]
port 167 nsew signal output
rlabel metal3 s 79200 132608 80000 132728 6 o_req_addr[14]
port 168 nsew signal output
rlabel metal3 s 79200 139408 80000 139528 6 o_req_addr[15]
port 169 nsew signal output
rlabel metal3 s 79200 36048 80000 36168 6 o_req_addr[1]
port 170 nsew signal output
rlabel metal3 s 79200 44208 80000 44328 6 o_req_addr[2]
port 171 nsew signal output
rlabel metal3 s 79200 52368 80000 52488 6 o_req_addr[3]
port 172 nsew signal output
rlabel metal3 s 79200 60528 80000 60648 6 o_req_addr[4]
port 173 nsew signal output
rlabel metal3 s 79200 68688 80000 68808 6 o_req_addr[5]
port 174 nsew signal output
rlabel metal3 s 79200 76848 80000 76968 6 o_req_addr[6]
port 175 nsew signal output
rlabel metal3 s 79200 85008 80000 85128 6 o_req_addr[7]
port 176 nsew signal output
rlabel metal3 s 79200 91808 80000 91928 6 o_req_addr[8]
port 177 nsew signal output
rlabel metal3 s 79200 98608 80000 98728 6 o_req_addr[9]
port 178 nsew signal output
rlabel metal3 s 79200 19048 80000 19168 6 o_req_ppl_submit
port 179 nsew signal output
rlabel metal3 s 79200 27888 80000 28008 6 sr_bus_addr[0]
port 180 nsew signal output
rlabel metal3 s 79200 106088 80000 106208 6 sr_bus_addr[10]
port 181 nsew signal output
rlabel metal3 s 79200 112888 80000 113008 6 sr_bus_addr[11]
port 182 nsew signal output
rlabel metal3 s 79200 119688 80000 119808 6 sr_bus_addr[12]
port 183 nsew signal output
rlabel metal3 s 79200 126488 80000 126608 6 sr_bus_addr[13]
port 184 nsew signal output
rlabel metal3 s 79200 133288 80000 133408 6 sr_bus_addr[14]
port 185 nsew signal output
rlabel metal3 s 79200 140088 80000 140208 6 sr_bus_addr[15]
port 186 nsew signal output
rlabel metal3 s 79200 36728 80000 36848 6 sr_bus_addr[1]
port 187 nsew signal output
rlabel metal3 s 79200 44888 80000 45008 6 sr_bus_addr[2]
port 188 nsew signal output
rlabel metal3 s 79200 53048 80000 53168 6 sr_bus_addr[3]
port 189 nsew signal output
rlabel metal3 s 79200 61208 80000 61328 6 sr_bus_addr[4]
port 190 nsew signal output
rlabel metal3 s 79200 69368 80000 69488 6 sr_bus_addr[5]
port 191 nsew signal output
rlabel metal3 s 79200 77528 80000 77648 6 sr_bus_addr[6]
port 192 nsew signal output
rlabel metal3 s 79200 85688 80000 85808 6 sr_bus_addr[7]
port 193 nsew signal output
rlabel metal3 s 79200 92488 80000 92608 6 sr_bus_addr[8]
port 194 nsew signal output
rlabel metal3 s 79200 99288 80000 99408 6 sr_bus_addr[9]
port 195 nsew signal output
rlabel metal3 s 79200 28568 80000 28688 6 sr_bus_data_o[0]
port 196 nsew signal output
rlabel metal3 s 79200 106768 80000 106888 6 sr_bus_data_o[10]
port 197 nsew signal output
rlabel metal3 s 79200 113568 80000 113688 6 sr_bus_data_o[11]
port 198 nsew signal output
rlabel metal3 s 79200 120368 80000 120488 6 sr_bus_data_o[12]
port 199 nsew signal output
rlabel metal3 s 79200 127168 80000 127288 6 sr_bus_data_o[13]
port 200 nsew signal output
rlabel metal3 s 79200 133968 80000 134088 6 sr_bus_data_o[14]
port 201 nsew signal output
rlabel metal3 s 79200 140768 80000 140888 6 sr_bus_data_o[15]
port 202 nsew signal output
rlabel metal3 s 79200 37408 80000 37528 6 sr_bus_data_o[1]
port 203 nsew signal output
rlabel metal3 s 79200 45568 80000 45688 6 sr_bus_data_o[2]
port 204 nsew signal output
rlabel metal3 s 79200 53728 80000 53848 6 sr_bus_data_o[3]
port 205 nsew signal output
rlabel metal3 s 79200 61888 80000 62008 6 sr_bus_data_o[4]
port 206 nsew signal output
rlabel metal3 s 79200 70048 80000 70168 6 sr_bus_data_o[5]
port 207 nsew signal output
rlabel metal3 s 79200 78208 80000 78328 6 sr_bus_data_o[6]
port 208 nsew signal output
rlabel metal3 s 79200 86368 80000 86488 6 sr_bus_data_o[7]
port 209 nsew signal output
rlabel metal3 s 79200 93168 80000 93288 6 sr_bus_data_o[8]
port 210 nsew signal output
rlabel metal3 s 79200 99968 80000 100088 6 sr_bus_data_o[9]
port 211 nsew signal output
rlabel metal3 s 79200 19728 80000 19848 6 sr_bus_we
port 212 nsew signal output
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 213 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 213 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 213 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 214 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 214 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 80000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 19040418
string GDS_FILE /home/piotro/caravel_user_project/openlane/core1/runs/22_12_31_15_08/results/signoff/core1.magic.gds
string GDS_START 1273108
<< end >>

