magic
tech sky130B
magscale 1 2
timestamp 1662802087
<< obsli1 >>
rect 1104 2159 198812 379729
<< obsm1 >>
rect 382 2128 199810 379760
<< obsm2 >>
rect 386 2139 199990 379749
<< metal3 >>
rect 199200 378088 200000 378208
rect 0 375096 800 375216
rect 199200 372240 200000 372360
rect 0 369248 800 369368
rect 199200 366392 200000 366512
rect 0 363400 800 363520
rect 199200 360544 200000 360664
rect 0 357552 800 357672
rect 199200 354696 200000 354816
rect 0 351704 800 351824
rect 199200 348848 200000 348968
rect 0 345856 800 345976
rect 199200 343000 200000 343120
rect 0 340008 800 340128
rect 199200 337152 200000 337272
rect 0 334160 800 334280
rect 199200 331304 200000 331424
rect 0 328312 800 328432
rect 199200 325456 200000 325576
rect 0 322464 800 322584
rect 199200 319608 200000 319728
rect 0 316616 800 316736
rect 199200 313760 200000 313880
rect 0 310768 800 310888
rect 199200 307912 200000 308032
rect 0 304920 800 305040
rect 199200 302064 200000 302184
rect 0 299072 800 299192
rect 199200 296216 200000 296336
rect 0 293224 800 293344
rect 199200 290368 200000 290488
rect 0 287376 800 287496
rect 199200 284520 200000 284640
rect 0 281528 800 281648
rect 199200 278672 200000 278792
rect 0 275680 800 275800
rect 199200 272824 200000 272944
rect 0 269832 800 269952
rect 199200 266976 200000 267096
rect 0 263984 800 264104
rect 199200 261128 200000 261248
rect 0 258136 800 258256
rect 199200 255280 200000 255400
rect 0 252288 800 252408
rect 199200 249432 200000 249552
rect 0 246440 800 246560
rect 199200 243584 200000 243704
rect 0 240592 800 240712
rect 199200 237736 200000 237856
rect 0 234744 800 234864
rect 199200 231888 200000 232008
rect 0 228896 800 229016
rect 199200 226040 200000 226160
rect 0 223048 800 223168
rect 199200 220192 200000 220312
rect 0 217200 800 217320
rect 199200 214344 200000 214464
rect 0 211352 800 211472
rect 199200 208496 200000 208616
rect 0 205504 800 205624
rect 199200 202648 200000 202768
rect 0 199656 800 199776
rect 199200 196800 200000 196920
rect 0 193808 800 193928
rect 199200 190952 200000 191072
rect 0 187960 800 188080
rect 199200 185104 200000 185224
rect 0 182112 800 182232
rect 199200 179256 200000 179376
rect 0 176264 800 176384
rect 199200 173408 200000 173528
rect 0 170416 800 170536
rect 199200 167560 200000 167680
rect 0 164568 800 164688
rect 199200 161712 200000 161832
rect 0 158720 800 158840
rect 199200 155864 200000 155984
rect 0 152872 800 152992
rect 199200 150016 200000 150136
rect 0 147024 800 147144
rect 199200 144168 200000 144288
rect 0 141176 800 141296
rect 199200 138320 200000 138440
rect 0 135328 800 135448
rect 199200 132472 200000 132592
rect 0 129480 800 129600
rect 199200 126624 200000 126744
rect 0 123632 800 123752
rect 199200 120776 200000 120896
rect 0 117784 800 117904
rect 199200 114928 200000 115048
rect 0 111936 800 112056
rect 199200 109080 200000 109200
rect 0 106088 800 106208
rect 199200 103232 200000 103352
rect 0 100240 800 100360
rect 199200 97384 200000 97504
rect 0 94392 800 94512
rect 199200 91536 200000 91656
rect 0 88544 800 88664
rect 199200 85688 200000 85808
rect 0 82696 800 82816
rect 199200 79840 200000 79960
rect 0 76848 800 76968
rect 199200 73992 200000 74112
rect 0 71000 800 71120
rect 199200 68144 200000 68264
rect 0 65152 800 65272
rect 199200 62296 200000 62416
rect 0 59304 800 59424
rect 199200 56448 200000 56568
rect 0 53456 800 53576
rect 199200 50600 200000 50720
rect 0 47608 800 47728
rect 199200 44752 200000 44872
rect 0 41760 800 41880
rect 199200 38904 200000 39024
rect 0 35912 800 36032
rect 199200 33056 200000 33176
rect 0 30064 800 30184
rect 199200 27208 200000 27328
rect 0 24216 800 24336
rect 199200 21360 200000 21480
rect 0 18368 800 18488
rect 199200 15512 200000 15632
rect 0 12520 800 12640
rect 199200 9664 200000 9784
rect 0 6672 800 6792
rect 199200 3816 200000 3936
<< obsm3 >>
rect 238 378288 199995 379745
rect 238 378008 199120 378288
rect 238 375296 199995 378008
rect 880 375016 199995 375296
rect 238 372440 199995 375016
rect 238 372160 199120 372440
rect 238 369448 199995 372160
rect 880 369168 199995 369448
rect 238 366592 199995 369168
rect 238 366312 199120 366592
rect 238 363600 199995 366312
rect 880 363320 199995 363600
rect 238 360744 199995 363320
rect 238 360464 199120 360744
rect 238 357752 199995 360464
rect 880 357472 199995 357752
rect 238 354896 199995 357472
rect 238 354616 199120 354896
rect 238 351904 199995 354616
rect 880 351624 199995 351904
rect 238 349048 199995 351624
rect 238 348768 199120 349048
rect 238 346056 199995 348768
rect 880 345776 199995 346056
rect 238 343200 199995 345776
rect 238 342920 199120 343200
rect 238 340208 199995 342920
rect 880 339928 199995 340208
rect 238 337352 199995 339928
rect 238 337072 199120 337352
rect 238 334360 199995 337072
rect 880 334080 199995 334360
rect 238 331504 199995 334080
rect 238 331224 199120 331504
rect 238 328512 199995 331224
rect 880 328232 199995 328512
rect 238 325656 199995 328232
rect 238 325376 199120 325656
rect 238 322664 199995 325376
rect 880 322384 199995 322664
rect 238 319808 199995 322384
rect 238 319528 199120 319808
rect 238 316816 199995 319528
rect 880 316536 199995 316816
rect 238 313960 199995 316536
rect 238 313680 199120 313960
rect 238 310968 199995 313680
rect 880 310688 199995 310968
rect 238 308112 199995 310688
rect 238 307832 199120 308112
rect 238 305120 199995 307832
rect 880 304840 199995 305120
rect 238 302264 199995 304840
rect 238 301984 199120 302264
rect 238 299272 199995 301984
rect 880 298992 199995 299272
rect 238 296416 199995 298992
rect 238 296136 199120 296416
rect 238 293424 199995 296136
rect 880 293144 199995 293424
rect 238 290568 199995 293144
rect 238 290288 199120 290568
rect 238 287576 199995 290288
rect 880 287296 199995 287576
rect 238 284720 199995 287296
rect 238 284440 199120 284720
rect 238 281728 199995 284440
rect 880 281448 199995 281728
rect 238 278872 199995 281448
rect 238 278592 199120 278872
rect 238 275880 199995 278592
rect 880 275600 199995 275880
rect 238 273024 199995 275600
rect 238 272744 199120 273024
rect 238 270032 199995 272744
rect 880 269752 199995 270032
rect 238 267176 199995 269752
rect 238 266896 199120 267176
rect 238 264184 199995 266896
rect 880 263904 199995 264184
rect 238 261328 199995 263904
rect 238 261048 199120 261328
rect 238 258336 199995 261048
rect 880 258056 199995 258336
rect 238 255480 199995 258056
rect 238 255200 199120 255480
rect 238 252488 199995 255200
rect 880 252208 199995 252488
rect 238 249632 199995 252208
rect 238 249352 199120 249632
rect 238 246640 199995 249352
rect 880 246360 199995 246640
rect 238 243784 199995 246360
rect 238 243504 199120 243784
rect 238 240792 199995 243504
rect 880 240512 199995 240792
rect 238 237936 199995 240512
rect 238 237656 199120 237936
rect 238 234944 199995 237656
rect 880 234664 199995 234944
rect 238 232088 199995 234664
rect 238 231808 199120 232088
rect 238 229096 199995 231808
rect 880 228816 199995 229096
rect 238 226240 199995 228816
rect 238 225960 199120 226240
rect 238 223248 199995 225960
rect 880 222968 199995 223248
rect 238 220392 199995 222968
rect 238 220112 199120 220392
rect 238 217400 199995 220112
rect 880 217120 199995 217400
rect 238 214544 199995 217120
rect 238 214264 199120 214544
rect 238 211552 199995 214264
rect 880 211272 199995 211552
rect 238 208696 199995 211272
rect 238 208416 199120 208696
rect 238 205704 199995 208416
rect 880 205424 199995 205704
rect 238 202848 199995 205424
rect 238 202568 199120 202848
rect 238 199856 199995 202568
rect 880 199576 199995 199856
rect 238 197000 199995 199576
rect 238 196720 199120 197000
rect 238 194008 199995 196720
rect 880 193728 199995 194008
rect 238 191152 199995 193728
rect 238 190872 199120 191152
rect 238 188160 199995 190872
rect 880 187880 199995 188160
rect 238 185304 199995 187880
rect 238 185024 199120 185304
rect 238 182312 199995 185024
rect 880 182032 199995 182312
rect 238 179456 199995 182032
rect 238 179176 199120 179456
rect 238 176464 199995 179176
rect 880 176184 199995 176464
rect 238 173608 199995 176184
rect 238 173328 199120 173608
rect 238 170616 199995 173328
rect 880 170336 199995 170616
rect 238 167760 199995 170336
rect 238 167480 199120 167760
rect 238 164768 199995 167480
rect 880 164488 199995 164768
rect 238 161912 199995 164488
rect 238 161632 199120 161912
rect 238 158920 199995 161632
rect 880 158640 199995 158920
rect 238 156064 199995 158640
rect 238 155784 199120 156064
rect 238 153072 199995 155784
rect 880 152792 199995 153072
rect 238 150216 199995 152792
rect 238 149936 199120 150216
rect 238 147224 199995 149936
rect 880 146944 199995 147224
rect 238 144368 199995 146944
rect 238 144088 199120 144368
rect 238 141376 199995 144088
rect 880 141096 199995 141376
rect 238 138520 199995 141096
rect 238 138240 199120 138520
rect 238 135528 199995 138240
rect 880 135248 199995 135528
rect 238 132672 199995 135248
rect 238 132392 199120 132672
rect 238 129680 199995 132392
rect 880 129400 199995 129680
rect 238 126824 199995 129400
rect 238 126544 199120 126824
rect 238 123832 199995 126544
rect 880 123552 199995 123832
rect 238 120976 199995 123552
rect 238 120696 199120 120976
rect 238 117984 199995 120696
rect 880 117704 199995 117984
rect 238 115128 199995 117704
rect 238 114848 199120 115128
rect 238 112136 199995 114848
rect 880 111856 199995 112136
rect 238 109280 199995 111856
rect 238 109000 199120 109280
rect 238 106288 199995 109000
rect 880 106008 199995 106288
rect 238 103432 199995 106008
rect 238 103152 199120 103432
rect 238 100440 199995 103152
rect 880 100160 199995 100440
rect 238 97584 199995 100160
rect 238 97304 199120 97584
rect 238 94592 199995 97304
rect 880 94312 199995 94592
rect 238 91736 199995 94312
rect 238 91456 199120 91736
rect 238 88744 199995 91456
rect 880 88464 199995 88744
rect 238 85888 199995 88464
rect 238 85608 199120 85888
rect 238 82896 199995 85608
rect 880 82616 199995 82896
rect 238 80040 199995 82616
rect 238 79760 199120 80040
rect 238 77048 199995 79760
rect 880 76768 199995 77048
rect 238 74192 199995 76768
rect 238 73912 199120 74192
rect 238 71200 199995 73912
rect 880 70920 199995 71200
rect 238 68344 199995 70920
rect 238 68064 199120 68344
rect 238 65352 199995 68064
rect 880 65072 199995 65352
rect 238 62496 199995 65072
rect 238 62216 199120 62496
rect 238 59504 199995 62216
rect 880 59224 199995 59504
rect 238 56648 199995 59224
rect 238 56368 199120 56648
rect 238 53656 199995 56368
rect 880 53376 199995 53656
rect 238 50800 199995 53376
rect 238 50520 199120 50800
rect 238 47808 199995 50520
rect 880 47528 199995 47808
rect 238 44952 199995 47528
rect 238 44672 199120 44952
rect 238 41960 199995 44672
rect 880 41680 199995 41960
rect 238 39104 199995 41680
rect 238 38824 199120 39104
rect 238 36112 199995 38824
rect 880 35832 199995 36112
rect 238 33256 199995 35832
rect 238 32976 199120 33256
rect 238 30264 199995 32976
rect 880 29984 199995 30264
rect 238 27408 199995 29984
rect 238 27128 199120 27408
rect 238 24416 199995 27128
rect 880 24136 199995 24416
rect 238 21560 199995 24136
rect 238 21280 199120 21560
rect 238 18568 199995 21280
rect 880 18288 199995 18568
rect 238 15712 199995 18288
rect 238 15432 199120 15712
rect 238 12720 199995 15432
rect 880 12440 199995 12720
rect 238 9864 199995 12440
rect 238 9584 199120 9864
rect 238 6872 199995 9584
rect 880 6592 199995 6872
rect 238 4016 199995 6592
rect 238 3736 199120 4016
rect 238 2143 199995 3736
<< metal4 >>
rect 4208 2128 4528 379760
rect 19568 2128 19888 379760
rect 34928 2128 35248 379760
rect 50288 2128 50608 379760
rect 65648 2128 65968 379760
rect 81008 2128 81328 379760
rect 96368 2128 96688 379760
rect 111728 2128 112048 379760
rect 127088 2128 127408 379760
rect 142448 2128 142768 379760
rect 157808 2128 158128 379760
rect 173168 2128 173488 379760
rect 188528 2128 188848 379760
<< obsm4 >>
rect 243 7923 4128 375597
rect 4608 7923 19488 375597
rect 19968 7923 34848 375597
rect 35328 7923 50208 375597
rect 50688 7923 65568 375597
rect 66048 7923 80928 375597
rect 81408 7923 96288 375597
rect 96768 7923 111648 375597
rect 112128 7923 127008 375597
rect 127488 7923 142368 375597
rect 142848 7923 157728 375597
rect 158208 7923 173088 375597
rect 173568 7923 188448 375597
rect 188928 7923 197189 375597
<< labels >>
rlabel metal3 s 199200 372240 200000 372360 6 i_clk
port 1 nsew signal input
rlabel metal3 s 199200 378088 200000 378208 6 i_rst
port 2 nsew signal input
rlabel metal3 s 199200 3816 200000 3936 6 mem_ack
port 3 nsew signal output
rlabel metal3 s 199200 9664 200000 9784 6 mem_addr[0]
port 4 nsew signal input
rlabel metal3 s 199200 68144 200000 68264 6 mem_addr[10]
port 5 nsew signal input
rlabel metal3 s 199200 73992 200000 74112 6 mem_addr[11]
port 6 nsew signal input
rlabel metal3 s 199200 79840 200000 79960 6 mem_addr[12]
port 7 nsew signal input
rlabel metal3 s 199200 85688 200000 85808 6 mem_addr[13]
port 8 nsew signal input
rlabel metal3 s 199200 91536 200000 91656 6 mem_addr[14]
port 9 nsew signal input
rlabel metal3 s 199200 97384 200000 97504 6 mem_addr[15]
port 10 nsew signal input
rlabel metal3 s 199200 103232 200000 103352 6 mem_addr[16]
port 11 nsew signal input
rlabel metal3 s 199200 109080 200000 109200 6 mem_addr[17]
port 12 nsew signal input
rlabel metal3 s 199200 114928 200000 115048 6 mem_addr[18]
port 13 nsew signal input
rlabel metal3 s 199200 120776 200000 120896 6 mem_addr[19]
port 14 nsew signal input
rlabel metal3 s 199200 15512 200000 15632 6 mem_addr[1]
port 15 nsew signal input
rlabel metal3 s 199200 126624 200000 126744 6 mem_addr[20]
port 16 nsew signal input
rlabel metal3 s 199200 132472 200000 132592 6 mem_addr[21]
port 17 nsew signal input
rlabel metal3 s 199200 138320 200000 138440 6 mem_addr[22]
port 18 nsew signal input
rlabel metal3 s 199200 144168 200000 144288 6 mem_addr[23]
port 19 nsew signal input
rlabel metal3 s 199200 21360 200000 21480 6 mem_addr[2]
port 20 nsew signal input
rlabel metal3 s 199200 27208 200000 27328 6 mem_addr[3]
port 21 nsew signal input
rlabel metal3 s 199200 33056 200000 33176 6 mem_addr[4]
port 22 nsew signal input
rlabel metal3 s 199200 38904 200000 39024 6 mem_addr[5]
port 23 nsew signal input
rlabel metal3 s 199200 44752 200000 44872 6 mem_addr[6]
port 24 nsew signal input
rlabel metal3 s 199200 50600 200000 50720 6 mem_addr[7]
port 25 nsew signal input
rlabel metal3 s 199200 56448 200000 56568 6 mem_addr[8]
port 26 nsew signal input
rlabel metal3 s 199200 62296 200000 62416 6 mem_addr[9]
port 27 nsew signal input
rlabel metal3 s 199200 150016 200000 150136 6 mem_cache_enable
port 28 nsew signal input
rlabel metal3 s 199200 155864 200000 155984 6 mem_exception
port 29 nsew signal output
rlabel metal3 s 199200 161712 200000 161832 6 mem_i_data[0]
port 30 nsew signal input
rlabel metal3 s 199200 220192 200000 220312 6 mem_i_data[10]
port 31 nsew signal input
rlabel metal3 s 199200 226040 200000 226160 6 mem_i_data[11]
port 32 nsew signal input
rlabel metal3 s 199200 231888 200000 232008 6 mem_i_data[12]
port 33 nsew signal input
rlabel metal3 s 199200 237736 200000 237856 6 mem_i_data[13]
port 34 nsew signal input
rlabel metal3 s 199200 243584 200000 243704 6 mem_i_data[14]
port 35 nsew signal input
rlabel metal3 s 199200 249432 200000 249552 6 mem_i_data[15]
port 36 nsew signal input
rlabel metal3 s 199200 167560 200000 167680 6 mem_i_data[1]
port 37 nsew signal input
rlabel metal3 s 199200 173408 200000 173528 6 mem_i_data[2]
port 38 nsew signal input
rlabel metal3 s 199200 179256 200000 179376 6 mem_i_data[3]
port 39 nsew signal input
rlabel metal3 s 199200 185104 200000 185224 6 mem_i_data[4]
port 40 nsew signal input
rlabel metal3 s 199200 190952 200000 191072 6 mem_i_data[5]
port 41 nsew signal input
rlabel metal3 s 199200 196800 200000 196920 6 mem_i_data[6]
port 42 nsew signal input
rlabel metal3 s 199200 202648 200000 202768 6 mem_i_data[7]
port 43 nsew signal input
rlabel metal3 s 199200 208496 200000 208616 6 mem_i_data[8]
port 44 nsew signal input
rlabel metal3 s 199200 214344 200000 214464 6 mem_i_data[9]
port 45 nsew signal input
rlabel metal3 s 199200 255280 200000 255400 6 mem_o_data[0]
port 46 nsew signal output
rlabel metal3 s 199200 313760 200000 313880 6 mem_o_data[10]
port 47 nsew signal output
rlabel metal3 s 199200 319608 200000 319728 6 mem_o_data[11]
port 48 nsew signal output
rlabel metal3 s 199200 325456 200000 325576 6 mem_o_data[12]
port 49 nsew signal output
rlabel metal3 s 199200 331304 200000 331424 6 mem_o_data[13]
port 50 nsew signal output
rlabel metal3 s 199200 337152 200000 337272 6 mem_o_data[14]
port 51 nsew signal output
rlabel metal3 s 199200 343000 200000 343120 6 mem_o_data[15]
port 52 nsew signal output
rlabel metal3 s 199200 261128 200000 261248 6 mem_o_data[1]
port 53 nsew signal output
rlabel metal3 s 199200 266976 200000 267096 6 mem_o_data[2]
port 54 nsew signal output
rlabel metal3 s 199200 272824 200000 272944 6 mem_o_data[3]
port 55 nsew signal output
rlabel metal3 s 199200 278672 200000 278792 6 mem_o_data[4]
port 56 nsew signal output
rlabel metal3 s 199200 284520 200000 284640 6 mem_o_data[5]
port 57 nsew signal output
rlabel metal3 s 199200 290368 200000 290488 6 mem_o_data[6]
port 58 nsew signal output
rlabel metal3 s 199200 296216 200000 296336 6 mem_o_data[7]
port 59 nsew signal output
rlabel metal3 s 199200 302064 200000 302184 6 mem_o_data[8]
port 60 nsew signal output
rlabel metal3 s 199200 307912 200000 308032 6 mem_o_data[9]
port 61 nsew signal output
rlabel metal3 s 199200 348848 200000 348968 6 mem_req
port 62 nsew signal input
rlabel metal3 s 199200 354696 200000 354816 6 mem_sel[0]
port 63 nsew signal input
rlabel metal3 s 199200 360544 200000 360664 6 mem_sel[1]
port 64 nsew signal input
rlabel metal3 s 199200 366392 200000 366512 6 mem_we
port 65 nsew signal input
rlabel metal4 s 4208 2128 4528 379760 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 379760 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 379760 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 379760 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 379760 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 379760 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 379760 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 379760 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 379760 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 379760 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 379760 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 379760 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 379760 6 vssd1
port 67 nsew ground bidirectional
rlabel metal3 s 0 6672 800 6792 6 wb_4_burst
port 68 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 wb_ack
port 69 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 wb_adr[0]
port 70 nsew signal output
rlabel metal3 s 0 76848 800 76968 6 wb_adr[10]
port 71 nsew signal output
rlabel metal3 s 0 82696 800 82816 6 wb_adr[11]
port 72 nsew signal output
rlabel metal3 s 0 88544 800 88664 6 wb_adr[12]
port 73 nsew signal output
rlabel metal3 s 0 94392 800 94512 6 wb_adr[13]
port 74 nsew signal output
rlabel metal3 s 0 100240 800 100360 6 wb_adr[14]
port 75 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 wb_adr[15]
port 76 nsew signal output
rlabel metal3 s 0 111936 800 112056 6 wb_adr[16]
port 77 nsew signal output
rlabel metal3 s 0 117784 800 117904 6 wb_adr[17]
port 78 nsew signal output
rlabel metal3 s 0 123632 800 123752 6 wb_adr[18]
port 79 nsew signal output
rlabel metal3 s 0 129480 800 129600 6 wb_adr[19]
port 80 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 wb_adr[1]
port 81 nsew signal output
rlabel metal3 s 0 135328 800 135448 6 wb_adr[20]
port 82 nsew signal output
rlabel metal3 s 0 141176 800 141296 6 wb_adr[21]
port 83 nsew signal output
rlabel metal3 s 0 147024 800 147144 6 wb_adr[22]
port 84 nsew signal output
rlabel metal3 s 0 152872 800 152992 6 wb_adr[23]
port 85 nsew signal output
rlabel metal3 s 0 30064 800 30184 6 wb_adr[2]
port 86 nsew signal output
rlabel metal3 s 0 35912 800 36032 6 wb_adr[3]
port 87 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 wb_adr[4]
port 88 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 wb_adr[5]
port 89 nsew signal output
rlabel metal3 s 0 53456 800 53576 6 wb_adr[6]
port 90 nsew signal output
rlabel metal3 s 0 59304 800 59424 6 wb_adr[7]
port 91 nsew signal output
rlabel metal3 s 0 65152 800 65272 6 wb_adr[8]
port 92 nsew signal output
rlabel metal3 s 0 71000 800 71120 6 wb_adr[9]
port 93 nsew signal output
rlabel metal3 s 0 158720 800 158840 6 wb_cyc
port 94 nsew signal output
rlabel metal3 s 0 164568 800 164688 6 wb_err
port 95 nsew signal input
rlabel metal3 s 0 170416 800 170536 6 wb_i_dat[0]
port 96 nsew signal input
rlabel metal3 s 0 228896 800 229016 6 wb_i_dat[10]
port 97 nsew signal input
rlabel metal3 s 0 234744 800 234864 6 wb_i_dat[11]
port 98 nsew signal input
rlabel metal3 s 0 240592 800 240712 6 wb_i_dat[12]
port 99 nsew signal input
rlabel metal3 s 0 246440 800 246560 6 wb_i_dat[13]
port 100 nsew signal input
rlabel metal3 s 0 252288 800 252408 6 wb_i_dat[14]
port 101 nsew signal input
rlabel metal3 s 0 258136 800 258256 6 wb_i_dat[15]
port 102 nsew signal input
rlabel metal3 s 0 176264 800 176384 6 wb_i_dat[1]
port 103 nsew signal input
rlabel metal3 s 0 182112 800 182232 6 wb_i_dat[2]
port 104 nsew signal input
rlabel metal3 s 0 187960 800 188080 6 wb_i_dat[3]
port 105 nsew signal input
rlabel metal3 s 0 193808 800 193928 6 wb_i_dat[4]
port 106 nsew signal input
rlabel metal3 s 0 199656 800 199776 6 wb_i_dat[5]
port 107 nsew signal input
rlabel metal3 s 0 205504 800 205624 6 wb_i_dat[6]
port 108 nsew signal input
rlabel metal3 s 0 211352 800 211472 6 wb_i_dat[7]
port 109 nsew signal input
rlabel metal3 s 0 217200 800 217320 6 wb_i_dat[8]
port 110 nsew signal input
rlabel metal3 s 0 223048 800 223168 6 wb_i_dat[9]
port 111 nsew signal input
rlabel metal3 s 0 263984 800 264104 6 wb_o_dat[0]
port 112 nsew signal output
rlabel metal3 s 0 322464 800 322584 6 wb_o_dat[10]
port 113 nsew signal output
rlabel metal3 s 0 328312 800 328432 6 wb_o_dat[11]
port 114 nsew signal output
rlabel metal3 s 0 334160 800 334280 6 wb_o_dat[12]
port 115 nsew signal output
rlabel metal3 s 0 340008 800 340128 6 wb_o_dat[13]
port 116 nsew signal output
rlabel metal3 s 0 345856 800 345976 6 wb_o_dat[14]
port 117 nsew signal output
rlabel metal3 s 0 351704 800 351824 6 wb_o_dat[15]
port 118 nsew signal output
rlabel metal3 s 0 269832 800 269952 6 wb_o_dat[1]
port 119 nsew signal output
rlabel metal3 s 0 275680 800 275800 6 wb_o_dat[2]
port 120 nsew signal output
rlabel metal3 s 0 281528 800 281648 6 wb_o_dat[3]
port 121 nsew signal output
rlabel metal3 s 0 287376 800 287496 6 wb_o_dat[4]
port 122 nsew signal output
rlabel metal3 s 0 293224 800 293344 6 wb_o_dat[5]
port 123 nsew signal output
rlabel metal3 s 0 299072 800 299192 6 wb_o_dat[6]
port 124 nsew signal output
rlabel metal3 s 0 304920 800 305040 6 wb_o_dat[7]
port 125 nsew signal output
rlabel metal3 s 0 310768 800 310888 6 wb_o_dat[8]
port 126 nsew signal output
rlabel metal3 s 0 316616 800 316736 6 wb_o_dat[9]
port 127 nsew signal output
rlabel metal3 s 0 357552 800 357672 6 wb_sel[0]
port 128 nsew signal output
rlabel metal3 s 0 363400 800 363520 6 wb_sel[1]
port 129 nsew signal output
rlabel metal3 s 0 369248 800 369368 6 wb_stb
port 130 nsew signal output
rlabel metal3 s 0 375096 800 375216 6 wb_we
port 131 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 200000 382000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 168207876
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/dcache/runs/22_09_10_10_56/results/signoff/dcache.magic.gds
string GDS_START 792240
<< end >>

