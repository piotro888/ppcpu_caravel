* NGSPICE file created from interconnect_inner.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

.subckt interconnect_inner c0_disable c0_i_core_int_sreg[0] c0_i_core_int_sreg[11]
+ c0_i_core_int_sreg[12] c0_i_core_int_sreg[13] c0_i_core_int_sreg[14] c0_i_core_int_sreg[15]
+ c0_i_core_int_sreg[1] c0_i_core_int_sreg[4] c0_i_core_int_sreg[5] c0_i_irq c0_i_mc_core_int
+ c0_i_mem_ack c0_i_mem_data[0] c0_i_mem_data[10] c0_i_mem_data[11] c0_i_mem_data[12]
+ c0_i_mem_data[13] c0_i_mem_data[14] c0_i_mem_data[15] c0_i_mem_data[1] c0_i_mem_data[2]
+ c0_i_mem_data[3] c0_i_mem_data[4] c0_i_mem_data[5] c0_i_mem_data[6] c0_i_mem_data[7]
+ c0_i_mem_data[8] c0_i_mem_data[9] c0_i_mem_exception c0_i_req_data[0] c0_i_req_data[10]
+ c0_i_req_data[11] c0_i_req_data[12] c0_i_req_data[13] c0_i_req_data[14] c0_i_req_data[15]
+ c0_i_req_data[16] c0_i_req_data[17] c0_i_req_data[18] c0_i_req_data[19] c0_i_req_data[1]
+ c0_i_req_data[20] c0_i_req_data[21] c0_i_req_data[22] c0_i_req_data[23] c0_i_req_data[24]
+ c0_i_req_data[25] c0_i_req_data[26] c0_i_req_data[27] c0_i_req_data[28] c0_i_req_data[29]
+ c0_i_req_data[2] c0_i_req_data[30] c0_i_req_data[31] c0_i_req_data[3] c0_i_req_data[4]
+ c0_i_req_data[5] c0_i_req_data[6] c0_i_req_data[7] c0_i_req_data[8] c0_i_req_data[9]
+ c0_i_req_data_valid c0_o_c_data_page c0_o_c_instr_long c0_o_c_instr_page c0_o_icache_flush
+ c0_o_instr_long_addr[0] c0_o_instr_long_addr[1] c0_o_instr_long_addr[2] c0_o_instr_long_addr[3]
+ c0_o_instr_long_addr[4] c0_o_instr_long_addr[5] c0_o_instr_long_addr[6] c0_o_instr_long_addr[7]
+ c0_o_mem_addr[0] c0_o_mem_addr[10] c0_o_mem_addr[11] c0_o_mem_addr[12] c0_o_mem_addr[13]
+ c0_o_mem_addr[14] c0_o_mem_addr[15] c0_o_mem_addr[1] c0_o_mem_addr[2] c0_o_mem_addr[3]
+ c0_o_mem_addr[4] c0_o_mem_addr[5] c0_o_mem_addr[6] c0_o_mem_addr[7] c0_o_mem_addr[8]
+ c0_o_mem_addr[9] c0_o_mem_data[0] c0_o_mem_data[10] c0_o_mem_data[11] c0_o_mem_data[12]
+ c0_o_mem_data[13] c0_o_mem_data[14] c0_o_mem_data[15] c0_o_mem_data[1] c0_o_mem_data[2]
+ c0_o_mem_data[3] c0_o_mem_data[4] c0_o_mem_data[5] c0_o_mem_data[6] c0_o_mem_data[7]
+ c0_o_mem_data[8] c0_o_mem_data[9] c0_o_mem_high_addr[0] c0_o_mem_high_addr[1] c0_o_mem_high_addr[2]
+ c0_o_mem_high_addr[3] c0_o_mem_high_addr[4] c0_o_mem_high_addr[5] c0_o_mem_high_addr[6]
+ c0_o_mem_high_addr[7] c0_o_mem_long_mode c0_o_mem_req c0_o_mem_sel[0] c0_o_mem_sel[1]
+ c0_o_mem_we c0_o_req_active c0_o_req_addr[0] c0_o_req_addr[10] c0_o_req_addr[11]
+ c0_o_req_addr[12] c0_o_req_addr[13] c0_o_req_addr[14] c0_o_req_addr[15] c0_o_req_addr[1]
+ c0_o_req_addr[2] c0_o_req_addr[3] c0_o_req_addr[4] c0_o_req_addr[5] c0_o_req_addr[6]
+ c0_o_req_addr[7] c0_o_req_addr[8] c0_o_req_addr[9] c0_o_req_ppl_submit c0_rst c0_sr_bus_addr[0]
+ c0_sr_bus_addr[10] c0_sr_bus_addr[11] c0_sr_bus_addr[12] c0_sr_bus_addr[13] c0_sr_bus_addr[14]
+ c0_sr_bus_addr[15] c0_sr_bus_addr[1] c0_sr_bus_addr[2] c0_sr_bus_addr[3] c0_sr_bus_addr[4]
+ c0_sr_bus_addr[5] c0_sr_bus_addr[6] c0_sr_bus_addr[7] c0_sr_bus_addr[8] c0_sr_bus_addr[9]
+ c0_sr_bus_data_o[0] c0_sr_bus_data_o[10] c0_sr_bus_data_o[11] c0_sr_bus_data_o[12]
+ c0_sr_bus_data_o[13] c0_sr_bus_data_o[14] c0_sr_bus_data_o[15] c0_sr_bus_data_o[1]
+ c0_sr_bus_data_o[2] c0_sr_bus_data_o[3] c0_sr_bus_data_o[4] c0_sr_bus_data_o[5]
+ c0_sr_bus_data_o[6] c0_sr_bus_data_o[7] c0_sr_bus_data_o[8] c0_sr_bus_data_o[9]
+ c0_sr_bus_we c1_dbg_pc[0] c1_dbg_pc[10] c1_dbg_pc[11] c1_dbg_pc[12] c1_dbg_pc[13]
+ c1_dbg_pc[14] c1_dbg_pc[15] c1_dbg_pc[1] c1_dbg_pc[2] c1_dbg_pc[3] c1_dbg_pc[4]
+ c1_dbg_pc[5] c1_dbg_pc[6] c1_dbg_pc[7] c1_dbg_pc[8] c1_dbg_pc[9] c1_dbg_r0[0] c1_dbg_r0[10]
+ c1_dbg_r0[11] c1_dbg_r0[12] c1_dbg_r0[13] c1_dbg_r0[14] c1_dbg_r0[15] c1_dbg_r0[1]
+ c1_dbg_r0[2] c1_dbg_r0[3] c1_dbg_r0[4] c1_dbg_r0[5] c1_dbg_r0[6] c1_dbg_r0[7] c1_dbg_r0[8]
+ c1_dbg_r0[9] c1_disable c1_i_core_int_sreg[0] c1_i_core_int_sreg[1] c1_i_core_int_sreg[6]
+ c1_i_core_int_sreg[7] c1_i_core_int_sreg[8] c1_i_core_int_sreg[9] c1_i_irq c1_i_mc_core_int
+ c1_i_mem_ack c1_i_mem_data[0] c1_i_mem_data[10] c1_i_mem_data[11] c1_i_mem_data[12]
+ c1_i_mem_data[13] c1_i_mem_data[14] c1_i_mem_data[15] c1_i_mem_data[1] c1_i_mem_data[2]
+ c1_i_mem_data[3] c1_i_mem_data[4] c1_i_mem_data[5] c1_i_mem_data[6] c1_i_mem_data[7]
+ c1_i_mem_data[8] c1_i_mem_data[9] c1_i_mem_exception c1_i_req_data[0] c1_i_req_data[10]
+ c1_i_req_data[11] c1_i_req_data[12] c1_i_req_data[13] c1_i_req_data[14] c1_i_req_data[15]
+ c1_i_req_data[16] c1_i_req_data[17] c1_i_req_data[18] c1_i_req_data[19] c1_i_req_data[1]
+ c1_i_req_data[20] c1_i_req_data[21] c1_i_req_data[22] c1_i_req_data[23] c1_i_req_data[24]
+ c1_i_req_data[25] c1_i_req_data[26] c1_i_req_data[27] c1_i_req_data[28] c1_i_req_data[29]
+ c1_i_req_data[2] c1_i_req_data[30] c1_i_req_data[31] c1_i_req_data[3] c1_i_req_data[4]
+ c1_i_req_data[5] c1_i_req_data[6] c1_i_req_data[7] c1_i_req_data[8] c1_i_req_data[9]
+ c1_i_req_data_valid c1_o_c_data_page c1_o_c_instr_long c1_o_c_instr_page c1_o_icache_flush
+ c1_o_instr_long_addr[0] c1_o_instr_long_addr[1] c1_o_instr_long_addr[2] c1_o_instr_long_addr[3]
+ c1_o_instr_long_addr[4] c1_o_instr_long_addr[5] c1_o_instr_long_addr[6] c1_o_instr_long_addr[7]
+ c1_o_mem_addr[0] c1_o_mem_addr[10] c1_o_mem_addr[11] c1_o_mem_addr[12] c1_o_mem_addr[13]
+ c1_o_mem_addr[14] c1_o_mem_addr[15] c1_o_mem_addr[1] c1_o_mem_addr[2] c1_o_mem_addr[3]
+ c1_o_mem_addr[4] c1_o_mem_addr[5] c1_o_mem_addr[6] c1_o_mem_addr[7] c1_o_mem_addr[8]
+ c1_o_mem_addr[9] c1_o_mem_data[0] c1_o_mem_data[10] c1_o_mem_data[11] c1_o_mem_data[12]
+ c1_o_mem_data[13] c1_o_mem_data[14] c1_o_mem_data[15] c1_o_mem_data[1] c1_o_mem_data[2]
+ c1_o_mem_data[3] c1_o_mem_data[4] c1_o_mem_data[5] c1_o_mem_data[6] c1_o_mem_data[7]
+ c1_o_mem_data[8] c1_o_mem_data[9] c1_o_mem_high_addr[0] c1_o_mem_high_addr[1] c1_o_mem_high_addr[2]
+ c1_o_mem_high_addr[3] c1_o_mem_high_addr[4] c1_o_mem_high_addr[5] c1_o_mem_high_addr[6]
+ c1_o_mem_high_addr[7] c1_o_mem_long_mode c1_o_mem_req c1_o_mem_sel[0] c1_o_mem_sel[1]
+ c1_o_mem_we c1_o_req_active c1_o_req_addr[0] c1_o_req_addr[10] c1_o_req_addr[11]
+ c1_o_req_addr[12] c1_o_req_addr[13] c1_o_req_addr[14] c1_o_req_addr[15] c1_o_req_addr[1]
+ c1_o_req_addr[2] c1_o_req_addr[3] c1_o_req_addr[4] c1_o_req_addr[5] c1_o_req_addr[6]
+ c1_o_req_addr[7] c1_o_req_addr[8] c1_o_req_addr[9] c1_o_req_ppl_submit c1_rst c1_sr_bus_addr[0]
+ c1_sr_bus_addr[10] c1_sr_bus_addr[11] c1_sr_bus_addr[12] c1_sr_bus_addr[13] c1_sr_bus_addr[14]
+ c1_sr_bus_addr[15] c1_sr_bus_addr[1] c1_sr_bus_addr[2] c1_sr_bus_addr[3] c1_sr_bus_addr[4]
+ c1_sr_bus_addr[5] c1_sr_bus_addr[6] c1_sr_bus_addr[7] c1_sr_bus_addr[8] c1_sr_bus_addr[9]
+ c1_sr_bus_data_o[0] c1_sr_bus_data_o[10] c1_sr_bus_data_o[11] c1_sr_bus_data_o[12]
+ c1_sr_bus_data_o[13] c1_sr_bus_data_o[14] c1_sr_bus_data_o[15] c1_sr_bus_data_o[1]
+ c1_sr_bus_data_o[2] c1_sr_bus_data_o[3] c1_sr_bus_data_o[4] c1_sr_bus_data_o[5]
+ c1_sr_bus_data_o[6] c1_sr_bus_data_o[7] c1_sr_bus_data_o[8] c1_sr_bus_data_o[9]
+ c1_sr_bus_we core_clock core_reset dcache_mem_ack dcache_mem_addr[0] dcache_mem_addr[10]
+ dcache_mem_addr[11] dcache_mem_addr[12] dcache_mem_addr[13] dcache_mem_addr[14]
+ dcache_mem_addr[15] dcache_mem_addr[16] dcache_mem_addr[17] dcache_mem_addr[18]
+ dcache_mem_addr[19] dcache_mem_addr[1] dcache_mem_addr[20] dcache_mem_addr[21] dcache_mem_addr[22]
+ dcache_mem_addr[23] dcache_mem_addr[2] dcache_mem_addr[3] dcache_mem_addr[4] dcache_mem_addr[5]
+ dcache_mem_addr[6] dcache_mem_addr[7] dcache_mem_addr[8] dcache_mem_addr[9] dcache_mem_cache_enable
+ dcache_mem_exception dcache_mem_i_data[0] dcache_mem_i_data[10] dcache_mem_i_data[11]
+ dcache_mem_i_data[12] dcache_mem_i_data[13] dcache_mem_i_data[14] dcache_mem_i_data[15]
+ dcache_mem_i_data[1] dcache_mem_i_data[2] dcache_mem_i_data[3] dcache_mem_i_data[4]
+ dcache_mem_i_data[5] dcache_mem_i_data[6] dcache_mem_i_data[7] dcache_mem_i_data[8]
+ dcache_mem_i_data[9] dcache_mem_o_data[0] dcache_mem_o_data[10] dcache_mem_o_data[11]
+ dcache_mem_o_data[12] dcache_mem_o_data[13] dcache_mem_o_data[14] dcache_mem_o_data[15]
+ dcache_mem_o_data[1] dcache_mem_o_data[2] dcache_mem_o_data[3] dcache_mem_o_data[4]
+ dcache_mem_o_data[5] dcache_mem_o_data[6] dcache_mem_o_data[7] dcache_mem_o_data[8]
+ dcache_mem_o_data[9] dcache_mem_req dcache_mem_sel[0] dcache_mem_sel[1] dcache_mem_we
+ dcache_rst dcache_wb_4_burst dcache_wb_ack dcache_wb_adr[0] dcache_wb_adr[10] dcache_wb_adr[11]
+ dcache_wb_adr[12] dcache_wb_adr[13] dcache_wb_adr[14] dcache_wb_adr[15] dcache_wb_adr[16]
+ dcache_wb_adr[17] dcache_wb_adr[18] dcache_wb_adr[19] dcache_wb_adr[1] dcache_wb_adr[20]
+ dcache_wb_adr[21] dcache_wb_adr[22] dcache_wb_adr[23] dcache_wb_adr[2] dcache_wb_adr[3]
+ dcache_wb_adr[4] dcache_wb_adr[5] dcache_wb_adr[6] dcache_wb_adr[7] dcache_wb_adr[8]
+ dcache_wb_adr[9] dcache_wb_cyc dcache_wb_err dcache_wb_i_dat[0] dcache_wb_i_dat[10]
+ dcache_wb_i_dat[11] dcache_wb_i_dat[12] dcache_wb_i_dat[13] dcache_wb_i_dat[14]
+ dcache_wb_i_dat[15] dcache_wb_i_dat[1] dcache_wb_i_dat[2] dcache_wb_i_dat[3] dcache_wb_i_dat[4]
+ dcache_wb_i_dat[5] dcache_wb_i_dat[6] dcache_wb_i_dat[7] dcache_wb_i_dat[8] dcache_wb_i_dat[9]
+ dcache_wb_o_dat[0] dcache_wb_o_dat[10] dcache_wb_o_dat[11] dcache_wb_o_dat[12] dcache_wb_o_dat[13]
+ dcache_wb_o_dat[14] dcache_wb_o_dat[15] dcache_wb_o_dat[1] dcache_wb_o_dat[2] dcache_wb_o_dat[3]
+ dcache_wb_o_dat[4] dcache_wb_o_dat[5] dcache_wb_o_dat[6] dcache_wb_o_dat[7] dcache_wb_o_dat[8]
+ dcache_wb_o_dat[9] dcache_wb_sel[0] dcache_wb_sel[1] dcache_wb_stb dcache_wb_we
+ ic0_mem_ack ic0_mem_addr[0] ic0_mem_addr[10] ic0_mem_addr[11] ic0_mem_addr[12] ic0_mem_addr[13]
+ ic0_mem_addr[14] ic0_mem_addr[15] ic0_mem_addr[1] ic0_mem_addr[2] ic0_mem_addr[3]
+ ic0_mem_addr[4] ic0_mem_addr[5] ic0_mem_addr[6] ic0_mem_addr[7] ic0_mem_addr[8]
+ ic0_mem_addr[9] ic0_mem_cache_flush ic0_mem_data[0] ic0_mem_data[10] ic0_mem_data[11]
+ ic0_mem_data[12] ic0_mem_data[13] ic0_mem_data[14] ic0_mem_data[15] ic0_mem_data[16]
+ ic0_mem_data[17] ic0_mem_data[18] ic0_mem_data[19] ic0_mem_data[1] ic0_mem_data[20]
+ ic0_mem_data[21] ic0_mem_data[22] ic0_mem_data[23] ic0_mem_data[24] ic0_mem_data[25]
+ ic0_mem_data[26] ic0_mem_data[27] ic0_mem_data[28] ic0_mem_data[29] ic0_mem_data[2]
+ ic0_mem_data[30] ic0_mem_data[31] ic0_mem_data[3] ic0_mem_data[4] ic0_mem_data[5]
+ ic0_mem_data[6] ic0_mem_data[7] ic0_mem_data[8] ic0_mem_data[9] ic0_mem_ppl_submit
+ ic0_mem_req ic0_rst ic0_wb_ack ic0_wb_adr[0] ic0_wb_adr[10] ic0_wb_adr[11] ic0_wb_adr[12]
+ ic0_wb_adr[13] ic0_wb_adr[14] ic0_wb_adr[15] ic0_wb_adr[1] ic0_wb_adr[2] ic0_wb_adr[3]
+ ic0_wb_adr[4] ic0_wb_adr[5] ic0_wb_adr[6] ic0_wb_adr[7] ic0_wb_adr[8] ic0_wb_adr[9]
+ ic0_wb_cyc ic0_wb_err ic0_wb_i_dat[0] ic0_wb_i_dat[10] ic0_wb_i_dat[11] ic0_wb_i_dat[12]
+ ic0_wb_i_dat[13] ic0_wb_i_dat[14] ic0_wb_i_dat[15] ic0_wb_i_dat[1] ic0_wb_i_dat[2]
+ ic0_wb_i_dat[3] ic0_wb_i_dat[4] ic0_wb_i_dat[5] ic0_wb_i_dat[6] ic0_wb_i_dat[7]
+ ic0_wb_i_dat[8] ic0_wb_i_dat[9] ic0_wb_sel[0] ic0_wb_sel[1] ic0_wb_stb ic0_wb_we
+ ic1_mem_ack ic1_mem_addr[0] ic1_mem_addr[10] ic1_mem_addr[11] ic1_mem_addr[12] ic1_mem_addr[13]
+ ic1_mem_addr[14] ic1_mem_addr[15] ic1_mem_addr[1] ic1_mem_addr[2] ic1_mem_addr[3]
+ ic1_mem_addr[4] ic1_mem_addr[5] ic1_mem_addr[6] ic1_mem_addr[7] ic1_mem_addr[8]
+ ic1_mem_addr[9] ic1_mem_cache_flush ic1_mem_data[0] ic1_mem_data[10] ic1_mem_data[11]
+ ic1_mem_data[12] ic1_mem_data[13] ic1_mem_data[14] ic1_mem_data[15] ic1_mem_data[16]
+ ic1_mem_data[17] ic1_mem_data[18] ic1_mem_data[19] ic1_mem_data[1] ic1_mem_data[20]
+ ic1_mem_data[21] ic1_mem_data[22] ic1_mem_data[23] ic1_mem_data[24] ic1_mem_data[25]
+ ic1_mem_data[26] ic1_mem_data[27] ic1_mem_data[28] ic1_mem_data[29] ic1_mem_data[2]
+ ic1_mem_data[30] ic1_mem_data[31] ic1_mem_data[3] ic1_mem_data[4] ic1_mem_data[5]
+ ic1_mem_data[6] ic1_mem_data[7] ic1_mem_data[8] ic1_mem_data[9] ic1_mem_ppl_submit
+ ic1_mem_req ic1_rst ic1_wb_ack ic1_wb_adr[0] ic1_wb_adr[10] ic1_wb_adr[11] ic1_wb_adr[12]
+ ic1_wb_adr[13] ic1_wb_adr[14] ic1_wb_adr[15] ic1_wb_adr[1] ic1_wb_adr[2] ic1_wb_adr[3]
+ ic1_wb_adr[4] ic1_wb_adr[5] ic1_wb_adr[6] ic1_wb_adr[7] ic1_wb_adr[8] ic1_wb_adr[9]
+ ic1_wb_cyc ic1_wb_err ic1_wb_i_dat[0] ic1_wb_i_dat[10] ic1_wb_i_dat[11] ic1_wb_i_dat[12]
+ ic1_wb_i_dat[13] ic1_wb_i_dat[14] ic1_wb_i_dat[15] ic1_wb_i_dat[1] ic1_wb_i_dat[2]
+ ic1_wb_i_dat[3] ic1_wb_i_dat[4] ic1_wb_i_dat[5] ic1_wb_i_dat[6] ic1_wb_i_dat[7]
+ ic1_wb_i_dat[8] ic1_wb_i_dat[9] ic1_wb_sel[0] ic1_wb_sel[1] ic1_wb_stb ic1_wb_we
+ inner_disable inner_embed_mode inner_ext_irq inner_wb_4_burst inner_wb_8_burst inner_wb_ack
+ inner_wb_adr[0] inner_wb_adr[10] inner_wb_adr[11] inner_wb_adr[12] inner_wb_adr[13]
+ inner_wb_adr[14] inner_wb_adr[15] inner_wb_adr[16] inner_wb_adr[17] inner_wb_adr[18]
+ inner_wb_adr[19] inner_wb_adr[1] inner_wb_adr[20] inner_wb_adr[21] inner_wb_adr[22]
+ inner_wb_adr[23] inner_wb_adr[2] inner_wb_adr[3] inner_wb_adr[4] inner_wb_adr[5]
+ inner_wb_adr[6] inner_wb_adr[7] inner_wb_adr[8] inner_wb_adr[9] inner_wb_cyc inner_wb_err
+ inner_wb_i_dat[0] inner_wb_i_dat[10] inner_wb_i_dat[11] inner_wb_i_dat[12] inner_wb_i_dat[13]
+ inner_wb_i_dat[14] inner_wb_i_dat[15] inner_wb_i_dat[1] inner_wb_i_dat[2] inner_wb_i_dat[3]
+ inner_wb_i_dat[4] inner_wb_i_dat[5] inner_wb_i_dat[6] inner_wb_i_dat[7] inner_wb_i_dat[8]
+ inner_wb_i_dat[9] inner_wb_o_dat[0] inner_wb_o_dat[10] inner_wb_o_dat[11] inner_wb_o_dat[12]
+ inner_wb_o_dat[13] inner_wb_o_dat[14] inner_wb_o_dat[15] inner_wb_o_dat[1] inner_wb_o_dat[2]
+ inner_wb_o_dat[3] inner_wb_o_dat[4] inner_wb_o_dat[5] inner_wb_o_dat[6] inner_wb_o_dat[7]
+ inner_wb_o_dat[8] inner_wb_o_dat[9] inner_wb_sel[0] inner_wb_sel[1] inner_wb_stb
+ inner_wb_we vccd1 vssd1 c1_i_core_int_sreg[11] c0_i_core_int_sreg[3] c0_i_core_int_sreg[2]
+ c1_i_core_int_sreg[10] c0_i_core_int_sreg[10] c0_i_core_int_sreg[9] c0_i_core_int_sreg[8]
+ c1_i_core_int_sreg[5] c0_i_core_int_sreg[7] c1_i_core_int_sreg[15] c1_i_core_int_sreg[4]
+ c1_i_core_int_sreg[3] c1_i_core_int_sreg[14] c0_i_core_int_sreg[6] c1_i_core_int_sreg[13]
+ c1_i_core_int_sreg[2] c1_i_core_int_sreg[12]
XANTENNA__3140__A1 net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_83_core_clock clknet_4_10__leaf_core_clock clknet_leaf_83_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3114__I _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3155_ net122 _0905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_78_1898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3086_ _0845_ net529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6286__CLK clknet_leaf_40_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _0487_ clknet_leaf_53_core_clock dmmu1.page_table\[4\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4640__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input108_I c1_o_c_instr_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6845_ _0418_ clknet_leaf_37_core_clock dmmu0.page_table\[1\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6776_ _0349_ clknet_leaf_104_core_clock dmmu0.long_off_reg\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3988_ net113 immu_1.high_addr_off\[3\] _1650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_50_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5727_ _2758_ _0378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_85_1814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6145__A1 _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5658_ dmmu0.long_off_reg\[3\] _1803_ _2716_ _2720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input73_I c0_o_req_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4609_ _2059_ _2090_ _2092_ immu_1.page_table\[13\]\[2\] _2095_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5589_ _1976_ _2396_ _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold340 dmmu0.page_table\[11\]\[12\] net1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_83_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold351 immu_1.page_table\[10\]\[6\] net1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold362 dmmu1.page_table\[5\]\[8\] net1096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold373 immu_0.page_table\[9\]\[4\] net1107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4459__A1 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5120__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3131__A1 _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6629__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_2038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_2704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_2250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_2715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5959__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_2014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__CLK clknet_leaf_104_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_1460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3895__S _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3198__A1 _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4395__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3737__A3 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7166__I net165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6070__I _2957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6136__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4698__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5895__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_2086 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_30_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_92_core_clock_I clknet_4_8__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4870__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4960_ _1817_ _2299_ _2302_ dmmu0.page_table\[7\]\[8\] _2311_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_1633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3911_ _1555_ _1557_ _1301_ _1575_ _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_50_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4891_ _2264_ _0036_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_28_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6630_ _0203_ clknet_leaf_29_core_clock dmmu0.page_table\[12\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6181__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3842_ _1433_ _1507_ _1508_ _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5178__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6561_ _0134_ clknet_leaf_20_core_clock immu_0.page_table\[5\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7076__I net360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3773_ _1410_ _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_15_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5512_ _2637_ _0284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6127__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6492_ _0065_ clknet_leaf_28_core_clock dmmu0.page_table\[14\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5443_ _2596_ _0256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput412 net412 c0_i_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput423 net423 c0_i_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput434 net434 c0_i_req_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5350__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5374_ _2453_ _2553_ _2555_ net953 _2558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput445 net445 c0_i_req_data[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput456 net456 c0_i_req_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7113_ net404 net581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3361__A1 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput467 net467 c1_i_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput478 net478 c1_i_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4325_ _1861_ _1911_ _1914_ immu_1.page_table\[2\]\[6\] _1921_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_1897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput489 net489 c1_i_req_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_61_1176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5638__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7044_ net280 net431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4256_ _1879_ _0595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3207_ _0883_ _0954_ _0940_ _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_78_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4187_ _1822_ _0583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input225_I dcache_mem_o_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3138_ _0887_ _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6921__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3069_ _0835_ net469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4613__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5810__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6828_ _0401_ clknet_leaf_43_core_clock dmmu1.page_table\[10\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4377__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6759_ _0332_ clknet_leaf_36_core_clock dmmu0.page_table\[5\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6301__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5877__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output444_I net444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold170 dmmu0.page_table\[0\]\[6\] net904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold181 immu_0.page_table\[4\]\[4\] net915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6451__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold192 dmmu1.page_table\[12\]\[6\] net926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4301__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_2209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3910__C _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_25_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6109__A1 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3591__A1 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5332__A2 _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_36_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4110_ _1301_ net325 _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_9_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5090_ _2387_ _0112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4041_ immu_0.page_table\[8\]\[9\] immu_0.page_table\[9\]\[9\] immu_0.page_table\[10\]\[9\]
+ immu_0.page_table\[11\]\[9\] _1463_ _1371_ _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3646__A2 net231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4843__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6045__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5992_ _2914_ _0487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4943_ _2301_ _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4932__B _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_23_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4874_ _1817_ _2242_ _2244_ dmmu0.page_table\[9\]\[8\] _2253_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6324__CLK clknet_leaf_70_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6613_ _0186_ clknet_leaf_12_core_clock immu_0.page_table\[1\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3825_ immu_0.page_table\[12\]\[3\] immu_0.page_table\[13\]\[3\] _1396_ _1492_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3267__C _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6544_ _0117_ clknet_leaf_22_core_clock immu_0.page_table\[7\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3756_ immu_0.page_table\[4\]\[1\] immu_0.page_table\[5\]\[1\] immu_0.page_table\[12\]\[1\]
+ immu_0.page_table\[13\]\[1\] _1424_ _1377_ _1425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_40_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5571__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6475_ _0048_ clknet_leaf_103_core_clock dmmu0.page_table\[8\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6474__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3687_ _1348_ net364 _1359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input175_I c1_o_req_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5426_ _2455_ _2582_ _2584_ dmmu0.page_table\[2\]\[3\] _2588_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3334__A1 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4531__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5357_ _2547_ _0219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_7_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input342_I ic1_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4308_ _1839_ _1891_ _1909_ _1910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5288_ _2507_ _0190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input36_I c0_o_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5087__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4239_ net208 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3637__A2 net260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3193__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_14__f_core_clock clknet_3_7_0_core_clock clknet_4_14__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_1323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5011__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_2002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6817__CLK clknet_leaf_67_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3573__A1 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output659_I net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3325__A1 net150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3420__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4825__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6027__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Left_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6347__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5250__A1 _1971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3100__I1 net27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3800__A2 _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3239__S1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6497__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3610_ inner_wb_arbiter.o_sel_sig _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_43_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5553__A2 _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _2083_ _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3541_ _1270_ net556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4761__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6260_ _0642_ clknet_leaf_90_core_clock immu_1.page_table\[4\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5305__A2 _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3472_ _0897_ _1210_ _1211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3316__A1 _1054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5211_ _1811_ _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4513__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6191_ _0573_ clknet_leaf_3_core_clock immu_0.page_table\[11\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5856__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5142_ _2418_ _0133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5069__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _2277_ _2367_ _2369_ net798 _2377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3619__A2 net266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4816__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4024_ net115 immu_1.high_addr_off\[5\] _1684_ _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_75_1654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3122__I _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ net199 _2889_ _2891_ dmmu1.page_table\[5\]\[11\] _2904_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4926_ _1837_ _2137_ _2286_ _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_34_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4857_ _2243_ _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_47_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input292_I ic0_mem_data[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_29_core_clock_I clknet_4_5__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3808_ _1446_ _1475_ _1476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4788_ _1817_ _2191_ _2193_ immu_0.page_table\[12\]\[8\] _2202_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6527_ _0100_ clknet_leaf_8_core_clock immu_0.page_table\[8\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_1723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3739_ net366 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_43_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6458_ _0031_ clknet_leaf_31_core_clock dmmu0.page_table\[9\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3307__A1 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5409_ _2577_ _0241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6389_ _0771_ clknet_leaf_79_core_clock immu_1.page_table\[10\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_2108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3166__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output407_I net407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_1727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5232__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3794__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4991__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5535__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7174__I net163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5299__A1 net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_2107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_31_core_clock_I clknet_4_7__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5471__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5223__A1 _1971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3085__I0 net125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5760_ _2777_ _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_57_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4711_ _1780_ _2154_ _2155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_29_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4982__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5691_ _2738_ _0362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4642_ _2063_ _2108_ _2110_ immu_1.page_table\[12\]\[4\] _2115_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4734__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4573_ _1870_ _2052_ _2054_ immu_1.page_table\[15\]\[10\] _2073_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6312_ _0694_ clknet_leaf_88_core_clock immu_1.page_table\[3\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3524_ _1261_ net533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_25_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6243_ _0625_ clknet_leaf_88_core_clock immu_1.page_table\[2\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3455_ _1193_ _1194_ _0906_ _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3117__I _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6174_ _3018_ _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3386_ net153 dmmu1.long_off_reg\[3\] _1127_ _1128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__6512__CLK clknet_leaf_6_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5125_ _2407_ _0127_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3560__I1 net56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input138_I c1_o_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3280__C _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5056_ _2366_ _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4265__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4007_ _1666_ _1667_ _1668_ _1669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_36_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6662__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input305_I ic0_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4017__A2 _1678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5958_ _2895_ _0472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3320__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4909_ _2276_ _0042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5889_ _1873_ _1874_ _2031_ _2855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_47_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5517__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6192__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3387__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput301 ic0_mem_data[31] net301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput312 ic0_wb_adr[12] net312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output524_I net524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput323 ic0_wb_adr[8] net323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xhold30 immu_0.page_table\[5\]\[4\] net764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput334 ic1_mem_data[12] net334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput345 ic1_mem_data[22] net345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold41 immu_1.page_table\[3\]\[6\] net775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput356 ic1_mem_data[3] net356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold52 dmmu0.page_table\[5\]\[2\] net786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput367 ic1_wb_adr[13] net367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold63 immu_0.page_table\[7\]\[3\] net797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput378 ic1_wb_adr[9] net378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold74 dmmu1.page_table\[15\]\[8\] net808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput389 inner_wb_i_dat[0] net389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xhold85 dmmu0.page_table\[9\]\[5\] net819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_76_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold96 dmmu1.page_table\[9\]\[7\] net830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_6_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_97_core_clock_I clknet_4_9__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_34_core_clock clknet_4_7__leaf_core_clock clknet_leaf_34_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3697__I _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3862__S1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_7_Left_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3519__A1 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4716__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5417__I _2581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_5 net373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3365__C _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6535__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3240_ _0985_ _0986_ _0907_ _0987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5141__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5692__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3542__I1 net43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3171_ _0889_ _0895_ _0914_ _0920_ _0921_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_59_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6685__CLK clknet_leaf_104_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_73_core_clock clknet_4_9__leaf_core_clock clknet_leaf_73_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_52_1768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5444__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6930_ _0503_ clknet_leaf_60_core_clock dmmu1.page_table\[3\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5995__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _0434_ clknet_leaf_50_core_clock dmmu1.page_table\[8\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7079__I net332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5812_ _2792_ _2802_ _2804_ dmmu1.page_table\[9\]\[6\] _2811_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6792_ _0365_ clknet_leaf_69_core_clock dmmu1.page_table\[13\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3302__S0 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3758__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5743_ _2768_ _0384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3853__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5674_ _2057_ _2726_ _2728_ net924 _2730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_1417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4625_ _2103_ _2090_ _2092_ immu_1.page_table\[13\]\[9\] _2104_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3275__C _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4556_ _2062_ _0712_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5380__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3507_ _0878_ _1239_ _1244_ _0862_ _1245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_64_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4487_ _1849_ _2014_ _2016_ net744 _2019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input255_I dcache_wb_cyc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6226_ _0608_ clknet_leaf_89_core_clock immu_1.page_table\[0\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3369__S0 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3438_ _0878_ _1175_ _1177_ _1178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4030__S1 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3533__I1 net39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6157_ _1860_ _3000_ _3002_ net1036 _3009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3369_ dmmu0.page_table\[8\]\[8\] dmmu0.page_table\[9\]\[8\] dmmu0.page_table\[10\]\[8\]
+ dmmu0.page_table\[11\]\[8\] _0865_ _0868_ _1111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5108_ _1790_ _2396_ _2397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6088_ _2968_ _0529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5039_ _2269_ _2352_ _2354_ net783 _2358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3997__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_2643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6408__CLK clknet_leaf_112_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_2654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5738__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_2075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4946__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output474_I net474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_2583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6163__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_2084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3221__I0 _0967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_2469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output641_I net641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5674__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput120 c1_o_mem_addr[11] net120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput131 c1_o_mem_addr[7] net131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput142 c1_o_mem_data[2] net142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput153 c1_o_mem_high_addr[3] net153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput164 c1_o_req_addr[0] net164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput175 c1_o_req_addr[5] net175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput186 c1_sr_bus_addr[14] net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4229__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5426__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput197 c1_sr_bus_data_o[0] net197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3421__S _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5977__A2 _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4401__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4410_ _1969_ _0659_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4165__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_2015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5390_ _2531_ _2552_ _2554_ net820 _2566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput605 net605 ic0_wb_i_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__5901__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput616 net616 ic0_wb_i_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_58_1944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput627 net627 ic1_mem_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_58_1955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput638 net638 ic1_mem_req vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4341_ _1846_ _1927_ _1929_ immu_1.page_table\[5\]\[1\] _1931_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6179__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput649 net649 ic1_wb_i_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_39_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7060_ net297 net448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5114__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4272_ _1887_ _0603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_39_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6011_ _1770_ _2923_ _2925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_78_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3223_ _0955_ _0961_ _0966_ _0970_ net522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_20_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3140__A2 net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3154_ _0897_ _0903_ _0904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3085_ net125 net20 _0842_ _0845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_1298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6913_ _0486_ clknet_leaf_55_core_clock dmmu1.page_table\[4\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4640__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6844_ _0417_ clknet_leaf_68_core_clock dmmu1.page_table\[9\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6700__CLK clknet_leaf_41_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6775_ _0348_ clknet_leaf_107_core_clock dmmu0.long_off_reg\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3987_ net113 immu_1.high_addr_off\[3\] _1649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_50_1763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5726_ _2049_ _2742_ _2744_ dmmu1.page_table\[12\]\[12\] _2758_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5657_ _2719_ _0347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6145__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input372_I ic1_wb_adr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6850__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4608_ _2094_ _0732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5588_ _2679_ _0318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input66_I c0_o_req_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold330 immu_0.page_table\[4\]\[3\] net1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3903__A1 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold341 dmmu0.page_table\[10\]\[1\] net1075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4539_ _2049_ _2032_ _2034_ net872 _2050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_1534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold352 immu_0.page_table\[13\]\[6\] net1086 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold363 dmmu0.page_table\[3\]\[1\] net1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold374 immu_0.page_table\[12\]\[4\] net1108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4459__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6209_ _0591_ clknet_leaf_80_core_clock immu_1.page_table\[9\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7189_ net393 net646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3131__A2 _0880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6230__CLK clknet_leaf_82_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_2705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_2716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5959__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3514__S0 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6380__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4919__B1 _2262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_2094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3198__A2 _0939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4395__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_2059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4147__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5344__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5895__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4698__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7182__I net401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_79_Left_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6723__CLK clknet_leaf_44_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4622__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3910_ _1378_ _1560_ _1574_ _1381_ _1575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_47_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4890_ _2258_ _2261_ _2263_ net756 _2264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_28_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3841_ _1474_ immu_1.page_table\[15\]\[3\] _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_15_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6873__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _0133_ clknet_leaf_9_core_clock immu_0.page_table\[5\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3772_ net366 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5583__B1 _2665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5511_ _2457_ _2630_ _2632_ dmmu0.page_table\[13\]\[4\] _2637_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6491_ _0064_ clknet_leaf_28_core_clock dmmu0.page_table\[14\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6127__A2 _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5442_ _1994_ _2581_ _2583_ net969 _2596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_1810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput413 net413 c0_i_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5373_ _2557_ _0225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput424 net424 c0_i_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput435 net435 c0_i_req_data[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput446 net446 c0_i_req_data[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_65_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput457 net457 c0_i_req_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7112_ net403 net580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4324_ _1920_ _0622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput468 net468 c1_i_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput479 net479 c1_i_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5638__A1 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7043_ net279 net430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4255_ _1824_ _1876_ _1878_ immu_1.page_table\[7\]\[0\] _1879_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6253__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3206_ _0951_ _0953_ _0878_ _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3744__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4186_ _1821_ _1791_ _1793_ immu_0.page_table\[11\]\[10\] _1822_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_1685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3137_ _0886_ _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_1549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input120_I c1_o_mem_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6063__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input218_I dcache_mem_o_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3068_ net216 _0831_ _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5810__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4613__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6827_ _0400_ clknet_leaf_45_core_clock dmmu1.page_table\[10\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3795__I _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4377__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_2081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6758_ _0331_ clknet_leaf_99_core_clock dmmu0.page_table\[6\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5709_ _2749_ _0369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6689_ _0262_ clknet_leaf_91_core_clock immu_1.high_addr_off\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5877__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_2076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold160 dmmu1.page_table\[11\]\[11\] net894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_63_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold171 dmmu1.page_table\[13\]\[8\] net905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold182 immu_1.page_table\[9\]\[7\] net916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold193 immu_1.page_table\[11\]\[0\] net927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_output437_I net437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4301__A1 net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6746__CLK clknet_leaf_32_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_36_core_clock_I clknet_4_7__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_5__f_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4065__B1 _1718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5652__I1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6896__CLK clknet_leaf_68_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7177__I net396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5404__I1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5565__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6109__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5317__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3591__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6276__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__S0 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_3__f_core_clock clknet_3_1_0_core_clock clknet_4_3__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4040_ immu_0.page_table\[12\]\[9\] immu_0.page_table\[13\]\[9\] immu_0.page_table\[14\]\[9\]
+ immu_0.page_table\[15\]\[9\] _1463_ _1371_ _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_40_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4843__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6045__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _2788_ _2907_ _2909_ dmmu1.page_table\[4\]\[4\] _2914_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_1680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ _2300_ _2298_ _2301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_34_1544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4873_ _2252_ _0030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4359__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6612_ _0185_ clknet_leaf_19_core_clock immu_0.page_table\[1\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3824_ immu_0.page_table\[8\]\[3\] immu_0.page_table\[9\]\[3\] immu_0.page_table\[10\]\[3\]
+ immu_0.page_table\[11\]\[3\] _1370_ _1372_ _1491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_28_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3755_ _1369_ _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_54_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6543_ _0116_ clknet_leaf_23_core_clock immu_0.page_table\[7\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6619__CLK clknet_leaf_24_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6474_ _0047_ clknet_leaf_13_core_clock dmmu0.page_table\[8\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3686_ _1356_ _1357_ _1358_ net683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_67_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Right_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5425_ _2587_ _0247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4531__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5356_ _2527_ _2536_ _2538_ net1105 _2547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input168_I c1_o_req_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6769__CLK clknet_leaf_99_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4307_ _1827_ net181 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
X_5287_ _1802_ _2502_ _2504_ immu_0.page_table\[0\]\[3\] _2507_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5087__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input335_I ic1_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4238_ _1865_ _0591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4295__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input29_I c0_o_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3193__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4169_ _1809_ _1792_ _1794_ immu_0.page_table\[11\]\[5\] _1810_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_65_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_21_Right_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_2110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5547__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5011__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_2003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6299__CLK clknet_leaf_85_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3573__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4770__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Right_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3474__B _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3956__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4286__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4825__A2 _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6027__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5786__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3649__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3261__A1 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4761__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3540_ net147 net42 _1267_ _1270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6911__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3471_ dmmu1.page_table\[4\]\[11\] dmmu1.page_table\[5\]\[11\] dmmu1.page_table\[6\]\[11\]
+ dmmu1.page_table\[7\]\[11\] _0888_ _0901_ _1210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5210_ _2460_ _0159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4513__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6190_ _3025_ _3026_ _3027_ _1895_ _0572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4513__B2 dmmu1.page_table\[14\]\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5710__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5141_ _2265_ _2414_ _2416_ immu_0.page_table\[5\]\[1\] _2418_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5069__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5072_ _2376_ _0105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4816__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4023_ _1651_ _1682_ _1683_ _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5974_ _2903_ _0480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_2075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_2086 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4925_ net195 net196 _1833_ _2286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__3252__A1 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6441__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4856_ _1980_ _2241_ _2243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_35_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3807_ immu_1.page_table\[4\]\[2\] immu_1.page_table\[5\]\[2\] immu_1.page_table\[6\]\[2\]
+ immu_1.page_table\[7\]\[2\] _1474_ _1469_ _1475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_7_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4787_ _2201_ _0804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input285_I ic0_mem_data[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6526_ _0099_ clknet_leaf_3_core_clock immu_0.page_table\[8\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3738_ _1407_ _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_30_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6457_ _0030_ clknet_leaf_25_core_clock dmmu0.page_table\[9\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3669_ _1302_ net375 _1345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_1009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3307__A2 _1049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5408_ immu_0.high_addr_off\[4\] _1806_ _2572_ _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3938__S0 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6388_ _0770_ clknet_leaf_74_core_clock immu_1.page_table\[10\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5339_ _2537_ _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_58_1831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3166__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6009__A1 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3491__A1 net51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_24_core_clock clknet_4_5__leaf_core_clock clknet_leaf_24_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_35_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5232__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4144__I _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4991__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6934__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4743__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5299__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7190__I net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_core_clock clknet_4_11__leaf_core_clock clknet_leaf_63_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6314__CLK clknet_leaf_70_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4259__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5471__A2 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6464__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4431__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4710_ net85 net84 _2154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4982__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5690_ _2103_ _2726_ _2728_ dmmu1.page_table\[13\]\[9\] _2738_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_84_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4641_ _2114_ _0745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4734__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4572_ _2072_ _0718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5931__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6311_ _0693_ clknet_leaf_88_core_clock immu_1.page_table\[3\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3523_ _1246_ _1260_ _0821_ _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6242_ _0624_ clknet_leaf_85_core_clock immu_1.page_table\[2\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_1610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3454_ dmmu1.page_table\[0\]\[10\] dmmu1.page_table\[1\]\[10\] dmmu1.page_table\[2\]\[10\]
+ dmmu1.page_table\[3\]\[10\] _0887_ _0909_ _1194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_21_880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6173_ dmmu1.long_off_reg\[1\] _1846_ _3016_ _3018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3385_ _1082_ _1125_ _1126_ _1127_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_42_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5124_ _2275_ _2398_ _2400_ immu_0.page_table\[6\]\[6\] _2407_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5055_ _1790_ _2259_ _2366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6807__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4006_ _1666_ _1667_ net2 _1668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4670__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input200_I c1_sr_bus_data_o[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6957__CLK clknet_leaf_62_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5957_ _2784_ _2890_ _2892_ dmmu1.page_table\[5\]\[2\] _2895_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3320__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4908_ _2275_ _2261_ _2263_ net906 _2276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5888_ _2854_ _0443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input96_I c0_sr_bus_data_o[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_33_Left_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4839_ _1812_ _2224_ _2226_ net1027 _2233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_51_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6509_ _0082_ clknet_leaf_4_core_clock immu_0.page_table\[10\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4489__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_1890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3387__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3244__S _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput302 ic0_mem_data[3] net302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_42_Left_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput313 ic0_wb_adr[13] net313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput324 ic0_wb_adr[9] net324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xhold20 dmmu0.page_table\[0\]\[9\] net754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput335 ic1_mem_data[13] net335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold31 immu_1.page_table\[15\]\[7\] net765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput346 ic1_mem_data[23] net346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold42 immu_1.page_table\[2\]\[8\] net776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput357 ic1_mem_data[4] net357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6487__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold53 dmmu0.page_table\[5\]\[9\] net787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_76_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold64 immu_0.page_table\[8\]\[7\] net798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput368 ic1_wb_adr[14] net368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5989__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput379 ic1_wb_cyc net379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xhold75 dmmu0.page_table\[6\]\[12\] net809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold86 dmmu0.page_table\[11\]\[10\] net820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold97 dmmu0.page_table\[15\]\[6\] net831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_19_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4075__S _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_51_Left_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4964__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7185__I net404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4716__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_6 net393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_2030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3662__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Left_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5141__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5692__A2 _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3170_ _0915_ _0917_ _0919_ _0920_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_52_1769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5444__A2 _2581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4652__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6860_ _0433_ clknet_leaf_49_core_clock dmmu1.page_table\[8\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_2012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5811_ _2810_ _0410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_2023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3207__A1 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6791_ _0364_ clknet_leaf_43_core_clock dmmu1.page_table\[13\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3302__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5742_ _2065_ _2760_ _2762_ dmmu1.page_table\[11\]\[5\] _2768_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_50_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6157__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5673_ _2729_ _0353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Right_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4624_ net209 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_13_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4183__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5380__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4555_ _2061_ _2053_ _2055_ immu_1.page_table\[15\]\[3\] _2062_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3128__I net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3506_ net18 _1241_ _1243_ _1244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_41_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3930__A2 _1582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4486_ _2018_ _0686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_1159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6225_ _0607_ clknet_leaf_81_core_clock immu_1.page_table\[0\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5132__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3437_ _0877_ _1176_ _1177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3369__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input150_I c1_o_mem_high_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input248_I dcache_wb_adr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3291__C _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3368_ dmmu0.page_table\[12\]\[8\] dmmu0.page_table\[13\]\[8\] dmmu0.page_table\[14\]\[8\]
+ dmmu0.page_table\[15\]\[8\] _0865_ _0868_ _1110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6156_ _3008_ _0557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3694__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5107_ _2172_ _2296_ _2396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3299_ _0897_ _1043_ _1044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6087_ _2794_ _2958_ _2960_ net838 _2968_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5038_ _2357_ _0090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input11_I c0_o_instr_long_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_2644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_2190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6989_ _0562_ clknet_leaf_73_core_clock immu_1.page_table\[8\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4946__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3749__A2 _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4422__I _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_2595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output467_I net467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3382__B1 _1119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output634_I net634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5674__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput110 c1_o_instr_long_addr[0] net110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3685__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput121 c1_o_mem_addr[12] net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput132 c1_o_mem_addr[8] net132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4882__B1 _2243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput143 c1_o_mem_data[3] net143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput154 c1_o_mem_high_addr[4] net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput165 c1_o_req_addr[10] net165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput176 c1_o_req_addr[6] net176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5426__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput187 c1_sr_bus_addr[15] net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput198 c1_sr_bus_data_o[10] net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3437__A1 _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_110_core_clock clknet_4_0__leaf_core_clock clknet_leaf_110_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3296__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6502__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3657__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_59_Right_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3376__C _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_43_core_clock_I clknet_4_12__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4165__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5362__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput606 net606 ic0_wb_i_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_61_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6652__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput617 net617 ic0_wb_i_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3912__A2 _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4340_ _1930_ _0628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput628 net628 ic1_mem_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput639 net639 ic1_rst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5114__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4271_ _1866_ _1876_ _1878_ immu_1.page_table\[7\]\[8\] _1887_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5163__I _2429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3222_ _0895_ _0969_ _0897_ _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6010_ _2923_ _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_78_1812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I c0_o_c_instr_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3676__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3220__S0 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3153_ dmmu1.page_table\[4\]\[0\] dmmu1.page_table\[5\]\[0\] dmmu1.page_table\[6\]\[0\]
+ dmmu1.page_table\[7\]\[0\] _0899_ _0902_ _0903_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3140__A3 net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3084_ _0844_ net518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4625__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6912_ _0485_ clknet_leaf_54_core_clock dmmu1.page_table\[4\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6843_ _0416_ clknet_leaf_66_core_clock dmmu1.page_table\[9\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4928__A1 net406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6774_ _0347_ clknet_leaf_106_core_clock dmmu0.long_off_reg\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_77_Right_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3986_ _1628_ _1647_ _1648_ net670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_1190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_1540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5725_ _2757_ _0377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__I net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input198_I c1_sr_bus_data_o[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5656_ dmmu0.long_off_reg\[2\] _1800_ _2716_ _2719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4607_ _2057_ _2090_ _2092_ net921 _2094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5587_ _2049_ _2663_ _2665_ dmmu1.page_table\[15\]\[12\] _2679_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input365_I ic1_wb_adr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold320 dmmu1.page_table\[1\]\[6\] net1054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold331 dmmu0.page_table\[7\]\[12\] net1065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4538_ net200 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xhold342 dmmu0.page_table\[12\]\[2\] net1076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold353 dmmu0.page_table\[14\]\[3\] net1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_7_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_70_2312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input59_I c0_o_req_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold364 dmmu1.page_table\[12\]\[5\] net1098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold375 immu_1.page_table\[9\]\[6\] net1109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5105__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4469_ _1860_ _1999_ _2001_ immu_1.page_table\[1\]\[6\] _2008_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_79_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6208_ _0590_ clknet_leaf_74_core_clock immu_1.page_table\[9\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3667__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7188_ net392 net645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4864__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6139_ _1895_ _2991_ _2997_ _2998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_5_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_2706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_2252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_2717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_2263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3514__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A1 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_2149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6525__CLK clknet_leaf_2_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4919__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5041__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output584_I net584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4395__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5592__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4152__I _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6675__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5344__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5895__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_1820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4607__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4083__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3830__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_28_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3840_ _1405_ immu_1.page_table\[14\]\[3\] _1507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5583__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3771_ _1439_ _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5510_ _2636_ _0283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6490_ _0063_ clknet_leaf_99_core_clock dmmu0.page_table\[7\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5441_ _2595_ _0255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput414 net414 c0_i_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5372_ _2451_ _2553_ _2555_ dmmu0.page_table\[11\]\[1\] _2557_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput425 net425 c0_i_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3897__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput436 net436 c0_i_req_data[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7111_ net402 net579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput447 net447 c0_i_req_data[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput458 net458 c0_i_req_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4323_ _1858_ _1911_ _1914_ net1010 _1920_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput469 net469 c1_i_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5099__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5638__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7042_ net278 net429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4254_ _1877_ _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3649__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3205_ dmmu0.page_table\[12\]\[2\] dmmu0.page_table\[13\]\[2\] dmmu0.page_table\[14\]\[2\]
+ dmmu0.page_table\[15\]\[2\] _0950_ _0952_ _0953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_38_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4185_ net93 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3744__S1 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5621__I _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6548__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3136_ net120 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_74_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6063__A2 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3067_ _0834_ net468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5271__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input113_I c1_o_instr_long_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5810__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6826_ _0399_ clknet_leaf_47_core_clock dmmu1.page_table\[10\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5023__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4377__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6757_ _0330_ clknet_leaf_13_core_clock dmmu0.page_table\[6\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3969_ net8 immu_0.high_addr_off\[3\] _1632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_45_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5708_ _2061_ _2743_ _2745_ net959 _2749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6688_ _0261_ clknet_leaf_92_core_clock immu_1.high_addr_off\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5639_ _2709_ _0339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5877__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_2055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3888__A1 net5 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3432__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold150 dmmu1.page_table\[11\]\[12\] net884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold161 immu_1.page_table\[4\]\[7\] net895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold172 dmmu0.page_table\[8\]\[6\] net906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold183 immu_0.page_table\[14\]\[10\] net917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold194 dmmu1.page_table\[3\]\[2\] net928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4837__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4301__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3499__S0 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3812__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5565__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3040__A2 net159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5317__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5868__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3879__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3974__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3670__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_1984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6045__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5990_ _2913_ _0486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6840__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4941_ _1769_ _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_8_1067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3829__C _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4872_ _1815_ _2242_ _2244_ dmmu0.page_table\[9\]\[7\] _2252_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6611_ _0184_ clknet_leaf_18_core_clock immu_0.page_table\[1\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6990__CLK clknet_leaf_104_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3823_ _1382_ _1489_ _1378_ _1490_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_74_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4006__B net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6542_ _0115_ clknet_leaf_27_core_clock immu_0.page_table\[7\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3754_ immu_0.page_table\[0\]\[1\] immu_0.page_table\[1\]\[1\] immu_0.page_table\[8\]\[1\]
+ immu_0.page_table\[9\]\[1\] _1396_ _1377_ _1423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_27_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6473_ _0046_ clknet_leaf_101_core_clock dmmu0.page_table\[8\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6220__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3685_ _1337_ net254 _1358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3564__C net533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5424_ _2453_ _2582_ _2584_ dmmu0.page_table\[2\]\[2\] _2587_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5355_ _2546_ _0218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4531__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3136__I net120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4306_ _1908_ _0616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5286_ _2506_ _0189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4237_ _1864_ _1841_ _1843_ net916 _1865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input230_I dcache_wb_4_burst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4295__A1 _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input328_I ic0_wb_stb vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4168_ _1808_ _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_1483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_14_core_clock clknet_4_6__leaf_core_clock clknet_leaf_14_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_69_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3119_ dmmu0.page_table\[4\]\[0\] dmmu0.page_table\[5\]\[0\] dmmu0.page_table\[6\]\[0\]
+ dmmu0.page_table\[7\]\[0\] _0865_ _0868_ _0869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_74_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4047__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4099_ _1535_ net275 _1757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5244__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3270__A2 _0858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6809_ _0382_ clknet_leaf_49_core_clock dmmu1.page_table\[11\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5547__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3405__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6713__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3956__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_53_core_clock clknet_4_15__leaf_core_clock clknet_leaf_53_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_24_1758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5483__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6027__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5786__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7188__I net392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6243__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_92_core_clock clknet_4_8__leaf_core_clock clknet_leaf_92_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4761__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3470_ _0915_ _1206_ _1208_ _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6393__CLK clknet_leaf_109_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_2072 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4513__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5710__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5140_ _2417_ _0132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5071_ _2275_ _2367_ _2369_ net1103 _2376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3324__I0 _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4022_ net114 immu_1.high_addr_off\[4\] _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4029__A1 _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5973_ _2851_ _2889_ _2891_ net1058 _2903_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4924_ _1788_ _2222_ _2284_ _2285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_48_937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5529__A1 _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4855_ _2241_ _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3806_ _1409_ _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_16_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4786_ _1815_ _2191_ _2193_ immu_0.page_table\[12\]\[7\] _2201_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6525_ _0098_ clknet_leaf_2_core_clock immu_0.page_table\[9\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3737_ net385 _1406_ net107 _1407_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_67_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input180_I c1_o_req_ppl_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3294__C _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input278_I ic0_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6456_ _0029_ clknet_leaf_15_core_clock dmmu0.page_table\[9\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3668_ _1342_ _1343_ _1344_ net679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_2014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5407_ _2576_ _0240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3938__S1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6387_ _0769_ clknet_leaf_74_core_clock immu_1.page_table\[10\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3599_ net213 _1219_ _1300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5338_ _2300_ _2535_ _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_60_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input41_I c0_o_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5269_ _1814_ _2486_ _2488_ immu_0.page_table\[1\]\[7\] _2496_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6009__A2 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5217__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6266__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output497_I net497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4991__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5457__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4743__A2 _2174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4160__I _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_48_core_clock_I clknet_4_13__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3554__I0 net139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4259__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6609__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5759__A1 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4431__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1072 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4982__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4640_ _2061_ _2108_ _2110_ immu_1.page_table\[12\]\[3\] _2114_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_37_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_100_core_clock_I clknet_4_3__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4734__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4571_ _1868_ _2053_ _2055_ net793 _2072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5931__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6310_ _0692_ clknet_leaf_85_core_clock immu_1.page_table\[3\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3522_ _0894_ _1250_ _1259_ _1260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_1909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6241_ _0623_ clknet_leaf_96_core_clock immu_1.page_table\[2\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3453_ dmmu1.page_table\[4\]\[10\] dmmu1.page_table\[5\]\[10\] dmmu1.page_table\[6\]\[10\]
+ dmmu1.page_table\[7\]\[10\] _0887_ _0909_ _1193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4042__S0 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ _3017_ _0564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3384_ net152 dmmu1.long_off_reg\[2\] _1126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3170__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5123_ _2406_ _0126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5054_ _2365_ _0098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6289__CLK clknet_leaf_100_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_50_core_clock_I clknet_4_13__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4005_ net9 immu_0.high_addr_off\[4\] _1667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4670__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4245__I net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5956_ _2894_ _0471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4907_ _1811_ _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_75_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5887_ _2049_ _2835_ _2837_ net938 _2854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input395_I inner_wb_i_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4838_ _2232_ _0015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input89_I c0_sr_bus_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4769_ _2190_ _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_43_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6508_ _0081_ clknet_leaf_4_core_clock immu_0.page_table\[10\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6439_ _0012_ clknet_leaf_17_core_clock dmmu0.page_table\[10\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4489__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3525__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3536__I0 net145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5686__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_2398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_4_core_clock clknet_4_1__leaf_core_clock clknet_leaf_4_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput303 ic0_mem_data[4] net303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold10 immu_1.page_table\[3\]\[2\] net744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput314 ic0_wb_adr[14] net314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput325 net735 net325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold21 dmmu0.page_table\[3\]\[5\] net755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5438__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold32 dmmu0.page_table\[6\]\[9\] net766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput336 ic1_mem_data[14] net336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput347 ic1_mem_data[24] net347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput358 ic1_mem_data[5] net358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold43 dmmu1.page_table\[9\]\[11\] net777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5989__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold54 dmmu0.page_table\[13\]\[6\] net788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput369 ic1_wb_adr[15] net369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold65 immu_1.page_table\[14\]\[5\] net799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold76 immu_1.page_table\[14\]\[8\] net810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold87 dmmu1.page_table\[0\]\[8\] net821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_58_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold98 dmmu0.page_table\[14\]\[2\] net832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_19_1624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6901__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_100_core_clock clknet_4_3__leaf_core_clock clknet_leaf_100_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4413__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5610__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4964__A2 _2298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4177__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4716__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5913__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_4_0_core_clock clknet_0_core_clock clknet_3_4_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_7 net393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3527__I0 net141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_2075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5141__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6431__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4652__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6581__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_2051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5810_ _2790_ _2802_ _2804_ net898 _2810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6790_ _0363_ clknet_leaf_42_core_clock dmmu1.page_table\[13\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_2046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5741_ _2767_ _0383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5672_ _2051_ _2726_ _2728_ net883 _2729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6157__A1 _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4623_ _2102_ _0739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4554_ _1851_ _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_5_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5380__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3391__A1 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3505_ _0875_ _1242_ _1243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_1788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4485_ _1846_ _2014_ _2016_ immu_1.page_table\[3\]\[1\] _2018_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6224_ _0606_ clknet_leaf_84_core_clock immu_1.page_table\[0\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3436_ dmmu0.page_table\[8\]\[10\] dmmu0.page_table\[9\]\[10\] dmmu0.page_table\[10\]\[10\]
+ dmmu0.page_table\[11\]\[10\] _0871_ _0866_ _1176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5132__A2 _2397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3143__A1 net124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6155_ _1857_ _3000_ _3002_ immu_1.page_table\[8\]\[5\] _3008_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3367_ _1094_ _1109_ net527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input143_I c1_o_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3694__A2 net233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5106_ _2395_ _0120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6086_ _2967_ _0528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6924__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3298_ dmmu1.page_table\[0\]\[5\] dmmu1.page_table\[1\]\[5\] dmmu1.page_table\[2\]\[5\]
+ dmmu1.page_table\[3\]\[5\] _0888_ _0910_ _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_5037_ _2267_ _2352_ _2354_ net763 _2357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_0_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input310_I ic0_wb_adr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_85_2770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_2781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_2792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6988_ _0561_ clknet_leaf_80_core_clock immu_1.page_table\[8\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4946__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5939_ _2847_ _2873_ _2875_ net826 _2884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_62_2077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6304__CLK clknet_leaf_82_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_79_2596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3382__A1 net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6454__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6171__I1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4331__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput100 c0_sr_bus_data_o[5] net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3054__I _0827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput111 c1_o_instr_long_addr[1] net111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput122 c1_o_mem_addr[13] net122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4882__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3685__A2 net254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput133 c1_o_mem_addr[9] net133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput144 c1_o_mem_data[4] net144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput155 c1_o_mem_high_addr[5] net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput166 c1_o_req_addr[11] net166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput177 c1_o_req_addr[7] net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput188 c1_sr_bus_addr[1] net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput199 c1_sr_bus_data_o[11] net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_32_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4937__A2 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3296__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6139__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5362__A2 _2535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput607 net607 ic0_wb_i_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput618 net618 ic0_wb_i_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput629 net629 ic1_mem_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_50_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ _1886_ _0602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5114__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6947__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3221_ _0967_ _0968_ _0912_ _0969_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_1182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3676__A2 net322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3220__S1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3152_ _0901_ _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_20_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3140__A4 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6075__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_0__f_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_3083_ net118 net13 _0842_ _0844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3428__A2 _1168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4625__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6911_ _0484_ clknet_leaf_56_core_clock dmmu1.page_table\[4\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6842_ _0415_ clknet_leaf_67_core_clock dmmu1.page_table\[9\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6327__CLK clknet_leaf_63_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_1828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6773_ _0346_ clknet_leaf_106_core_clock dmmu0.long_off_reg\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3985_ _1535_ net241 _1648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5724_ _2047_ _2742_ _2744_ net770 _2757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5655_ _2718_ _0346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3139__I _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6477__CLK clknet_leaf_105_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4606_ _2093_ _0731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5586_ _2678_ _0317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3364__A1 net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold310 immu_1.page_table\[9\]\[1\] net1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold321 immu_1.page_table\[5\]\[8\] net1055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4561__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4537_ _2048_ _0707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold332 immu_1.page_table\[6\]\[2\] net1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold343 dmmu0.page_table\[13\]\[8\] net1077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input260_I dcache_wb_o_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold354 dmmu1.page_table\[11\]\[3\] net1088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5105__A2 _2381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input358_I ic1_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold365 immu_0.page_table\[3\]\[7\] net1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4468_ _2007_ _0679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4313__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6207_ _0589_ clknet_leaf_74_core_clock immu_1.page_table\[9\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3419_ dmmu1.page_table\[12\]\[9\] dmmu1.page_table\[13\]\[9\] dmmu1.page_table\[14\]\[9\]
+ dmmu1.page_table\[15\]\[9\] _0887_ _0900_ _1160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7187_ net391 net644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4399_ _1855_ _1957_ _1959_ net760 _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4864__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3667__A2 net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6138_ _2994_ _0809_ _0810_ _2997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_5_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _1828_ _1891_ _2030_ _2957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__3602__I _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_2707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_2253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_2718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A2 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_2030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3758__B _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4919__A2 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5041__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5592__A2 _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5465__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5344__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3355__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4552__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3107__A1 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_2023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_1810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_2078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6057__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4607__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5804__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4083__A2 net245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5280__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_1625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3830__A2 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_28_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3770_ _1416_ _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_32_1473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5583__A2 _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ _2531_ _2581_ _2583_ dmmu0.page_table\[2\]\[10\] _2595_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5371_ _2556_ _0224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput415 net415 c0_i_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput426 net426 c0_i_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7110_ net401 net578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput437 net437 c0_i_req_data[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput448 net448 c0_i_req_data[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4322_ _1919_ _0621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput459 net459 c0_i_req_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5099__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7041_ net308 net459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4253_ _1771_ _1875_ _1877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3649__A2 net316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3204_ _0867_ _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4184_ _1820_ _0582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3135_ _0882_ _0883_ _0884_ _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_78_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3066_ net215 _0831_ _0834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_56_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5271__A1 net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input106_I c1_o_c_data_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6825_ _0398_ clknet_leaf_51_core_clock dmmu1.page_table\[10\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5023__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3968_ _1581_ _1629_ _1630_ _1631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6756_ _0329_ clknet_leaf_13_core_clock dmmu0.page_table\[6\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3585__A1 net229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5707_ _2748_ _0368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4782__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6687_ _0260_ clknet_leaf_91_core_clock immu_1.high_addr_off\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_2500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3899_ _1463_ immu_0.page_table\[13\]\[5\] _1564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_2511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5638_ _1814_ _2699_ _2701_ net791 _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input71_I c0_o_req_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3337__A1 net151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_2023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5569_ _2061_ _2664_ _2666_ dmmu1.page_table\[15\]\[3\] _2670_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3432__S1 _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold140 immu_1.page_table\[11\]\[7\] net874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold151 dmmu0.page_table\[15\]\[2\] net885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold162 immu_0.page_table\[15\]\[4\] net896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_43_core_clock clknet_4_12__leaf_core_clock clknet_leaf_43_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold173 immu_1.page_table\[14\]\[10\] net907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold184 immu_0.page_table\[3\]\[10\] net918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold195 dmmu1.page_table\[0\]\[6\] net929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_79_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3533__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4837__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_2103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3499__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6642__CLK clknet_leaf_32_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5565__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6792__CLK clknet_leaf_69_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3120__S0 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_82_core_clock clknet_4_10__leaf_core_clock clknet_leaf_82_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_49_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5317__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_105_core_clock_I clknet_4_2__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4525__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_36_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3187__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5253__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_55_core_clock_I clknet_4_15__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4940_ _2298_ _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_73_1584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ _2251_ _0029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5005__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6610_ _0183_ clknet_leaf_17_core_clock immu_0.page_table\[1\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3822_ _1486_ _1488_ _1366_ _1489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3567__A1 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6541_ _0114_ clknet_leaf_21_core_clock immu_0.page_table\[7\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3753_ icache_arbiter.o_sel_sig _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_42_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6472_ _0045_ clknet_leaf_12_core_clock dmmu0.page_table\[8\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3684_ _1350_ net324 _1326_ _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3319__A1 _1052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5423_ _2586_ _0246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5354_ _2463_ _2536_ _2538_ net1067 _2546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_80_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4305_ net198 _1893_ _1896_ immu_1.page_table\[0\]\[10\] _1908_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3861__B _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5285_ _1799_ _2502_ _2504_ immu_0.page_table\[0\]\[2\] _2506_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3178__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4236_ _1863_ _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4295__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4248__I net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3152__I _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6665__CLK clknet_leaf_110_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4167_ net100 _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_input223_I dcache_mem_o_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3118_ _0867_ _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4098_ _1350_ net329 _1360_ _1756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5244__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3049_ net222 _0822_ _0825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_2101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6808_ _0381_ clknet_leaf_49_core_clock dmmu1.page_table\[11\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5547__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_2055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4755__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _0312_ clknet_leaf_46_core_clock dmmu1.page_table\[15\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_1477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3405__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5180__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output442_I net442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3730__A1 _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4286__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5483__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5786__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3797__A1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3341__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4994__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_1719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4621__I net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_core_clock core_clock clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_52_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5710__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6688__CLK clknet_leaf_92_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5070_ _2375_ _0104_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4021_ net114 immu_1.high_addr_off\[4\] _1682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3324__I1 _1065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5226__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3700__I _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5972_ _2902_ _0479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3332__S0 _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4923_ _1974_ _1782_ _1784_ _2284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_74_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4854_ _1977_ _2240_ _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_12_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3805_ _1408_ _1472_ _1434_ _1473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_27_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4785_ _2200_ _0803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3736_ net108 _1406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6524_ _0097_ clknet_leaf_5_core_clock immu_0.page_table\[9\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3667_ _1337_ net250 _1344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3147__I _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6455_ _0028_ clknet_leaf_25_core_clock dmmu0.page_table\[9\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input173_I c1_o_req_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5406_ immu_0.high_addr_off\[3\] _1803_ _2572_ _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6386_ _0768_ clknet_leaf_79_core_clock immu_1.page_table\[10\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3598_ _1299_ net417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5337_ _2535_ _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3083__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input340_I ic1_mem_data[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5268_ _2495_ _0182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input34_I c0_o_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4219_ net203 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5199_ _1799_ _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6009__A3 _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5217__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3323__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4976__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4728__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6830__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3554__I1 net34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4259__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6980__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6210__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__A2 _2137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3314__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4431__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6360__CLK clknet_leaf_63_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3676__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3395__C _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5392__B1 _2554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4570_ _2071_ _0717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5931__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3521_ net123 _1253_ _1258_ _0934_ _1259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_53_996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6240_ _0622_ clknet_leaf_89_core_clock immu_1.page_table\[2\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3452_ _1187_ _1190_ _1192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4042__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6171_ dmmu1.long_off_reg\[0\] _1824_ _3016_ _3017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3383_ net152 dmmu1.long_off_reg\[2\] _1125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5122_ _2273_ _2398_ _2400_ net1035 _2406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5447__A1 net325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5053_ _2332_ _2351_ _2353_ net887 _2365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4004_ _1631_ _1632_ _1665_ _1666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_79_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4670__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3430__I _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4958__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6703__CLK clknet_leaf_41_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5955_ _2782_ _2890_ _2892_ net823 _2894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ _2274_ _0041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5886_ _2853_ _0442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4837_ _1809_ _2224_ _2226_ net1007 _2232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input290_I ic0_mem_data[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4186__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input388_I inner_wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6853__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4768_ _1790_ _2189_ _2190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_44_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_1403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6507_ _0080_ clknet_leaf_2_core_clock immu_0.page_table\[10\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3719_ _1370_ immu_0.page_table\[2\]\[0\] _1389_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_70_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4699_ _2148_ _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_1556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6438_ _0011_ clknet_leaf_26_core_clock dmmu0.page_table\[10\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4489__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5686__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3536__I1 net40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6369_ _0751_ clknet_leaf_78_core_clock immu_1.page_table\[12\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_2399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput304 ic0_mem_data[5] net304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_1155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3792__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput315 ic0_wb_adr[15] net315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold11 dmmu1.page_table\[6\]\[3\] net745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput326 ic0_wb_sel[0] net326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5438__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold22 dmmu0.page_table\[8\]\[0\] net756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold33 dmmu0.page_table\[9\]\[6\] net767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput337 ic1_mem_data[15] net337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput348 ic1_mem_data[25] net348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold44 dmmu1.page_table\[1\]\[9\] net778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold55 immu_0.page_table\[9\]\[8\] net789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput359 ic1_mem_data[6] net359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5989__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold66 immu_0.page_table\[9\]\[9\] net800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4110__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold77 dmmu1.page_table\[12\]\[9\] net811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold88 immu_0.page_table\[10\]\[3\] net822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold99 dmmu0.page_table\[3\]\[2\] net833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_output405_I net405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_2015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_4_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6383__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5610__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4413__A2 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5461__I1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4177__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_8 net393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5126__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_2070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4101__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6726__CLK clknet_leaf_40_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4652__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5740_ _2063_ _2760_ _2762_ dmmu1.page_table\[11\]\[4\] _2767_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_6_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3463__I0 _1186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6157__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5671_ _2727_ _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_72_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4622_ _2101_ _2090_ _2092_ net1093 _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4553_ _2060_ _0711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_83_1734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3504_ dmmu0.page_table\[12\]\[12\] dmmu0.page_table\[13\]\[12\] dmmu0.page_table\[14\]\[12\]
+ dmmu0.page_table\[15\]\[12\] _0863_ net16 _1242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4484_ _2017_ _0685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5668__A1 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6223_ _0605_ clknet_leaf_94_core_clock immu_1.page_table\[7\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3435_ _0875_ _1174_ _1175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6256__CLK clknet_leaf_95_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6154_ _3007_ _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3774__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3366_ _0860_ _1103_ _1108_ _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_42_1497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5105_ _2332_ _2381_ _2383_ net977 _2395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6085_ _2792_ _2958_ _2960_ net1054 _2967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3297_ _0907_ _1041_ _1042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_77_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6093__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input136_I c1_o_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5036_ _2356_ _0089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__A1 _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3160__I _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_2771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input303_I ic0_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6987_ _0560_ clknet_leaf_79_core_clock immu_1.page_table\[8\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_66_2192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_2067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5938_ _2883_ _0464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_62_2078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5869_ _2843_ _0435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5356__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3906__A1 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3536__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3382__A2 net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4331__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput101 c0_sr_bus_data_o[6] net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput112 c1_o_instr_long_addr[2] net112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output522_I net522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput123 c1_o_mem_addr[14] net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4882__A2 _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput134 c1_o_mem_data[0] net134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3271__S _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput145 c1_o_mem_data[5] net145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput156 c1_o_mem_high_addr[6] net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_51_1760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput167 c1_o_req_addr[12] net167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput178 c1_o_req_addr[8] net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput189 c1_sr_bus_addr[2] net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_32_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3070__A1 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6279__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput608 net608 ic0_wb_i_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput619 net619 ic0_wb_i_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_58_1947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3220_ dmmu1.page_table\[12\]\[2\] dmmu1.page_table\[13\]\[2\] dmmu1.page_table\[14\]\[2\]
+ dmmu1.page_table\[15\]\[2\] _0889_ _0931_ _0968_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3756__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3151_ _0900_ _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_59_1202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6075__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3082_ _0843_ net562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4625__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5822__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6910_ _0483_ clknet_leaf_55_core_clock dmmu1.page_table\[4\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_112_core_clock_I clknet_4_0__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6841_ _0414_ clknet_leaf_43_core_clock dmmu1.page_table\[9\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4389__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6772_ _0345_ clknet_leaf_106_core_clock dmmu0.long_off_reg\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3984_ _1636_ _1646_ _1360_ _1647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5723_ _2756_ _0376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_85_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5654_ dmmu0.long_off_reg\[1\] _1797_ _2716_ _2718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5889__A1 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4605_ _2051_ _2090_ _2092_ net1040 _2093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5585_ _2047_ _2663_ _2665_ net974 _2678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold300 dmmu1.page_table\[8\]\[4\] net1034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4561__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold311 dmmu1.page_table\[9\]\[10\] net1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4536_ _2047_ _2032_ _2034_ dmmu1.page_table\[14\]\[11\] _2048_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold322 dmmu0.page_table\[5\]\[11\] net1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_leaf_62_core_clock_I clknet_4_14__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_33_core_clock clknet_4_7__leaf_core_clock clknet_leaf_33_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold333 dmmu0.page_table\[15\]\[7\] net1067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold344 dmmu0.page_table\[6\]\[0\] net1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_83_1597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold355 dmmu1.page_table\[10\]\[3\] net1089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold366 dmmu1.page_table\[0\]\[2\] net1100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4467_ _1857_ _1999_ _2001_ immu_1.page_table\[1\]\[5\] _2007_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3155__I net122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input253_I dcache_wb_adr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4313__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6206_ _0588_ clknet_leaf_80_core_clock immu_1.page_table\[9\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_1862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3747__S0 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3418_ _0894_ _1158_ _1159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_2014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4398_ _1963_ _0653_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7186_ net390 net643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4864__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6137_ _2996_ _0550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3349_ _0915_ _1086_ _1091_ _0894_ _1092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3091__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ _2956_ _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_83_2708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5664__I1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_2719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ _2275_ _2337_ _2339_ immu_0.page_table\[10\]\[6\] _2346_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_68_2265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_2129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5577__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5041__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_2007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_72_core_clock clknet_4_9__leaf_core_clock clknet_leaf_72_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_63_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Left_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4552__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6571__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_2051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_1800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3107__A2 net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6057__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5804__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4607__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_48_Left_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_1880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3130__I2 _0873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3291__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4624__I net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5656__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4240__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3684__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_57_Left_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6914__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5370_ _2444_ _2553_ _2555_ dmmu0.page_table\[11\]\[0\] _2556_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5740__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3977__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput405 net405 c0_disable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput416 net416 c0_i_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput427 net427 c0_i_mem_exception vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput438 net438 c0_i_req_data[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4321_ _1855_ _1911_ _1914_ immu_1.page_table\[2\]\[4\] _1919_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput449 net449 c0_i_req_data[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5099__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4252_ _1875_ _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7040_ net307 net458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3203_ dmmu0.page_table\[4\]\[2\] dmmu0.page_table\[5\]\[2\] dmmu0.page_table\[6\]\[2\]
+ dmmu0.page_table\[7\]\[2\] _0950_ _0948_ _0951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_43_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4183_ _1819_ _1792_ _1794_ immu_0.page_table\[11\]\[9\] _1820_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3134_ _0821_ _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_39_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_66_Left_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3065_ _0833_ net482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5271__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6444__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6824_ _0397_ clknet_leaf_50_core_clock dmmu1.page_table\[10\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5023__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6755_ _0328_ clknet_leaf_14_core_clock dmmu0.page_table\[6\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3967_ net7 immu_0.high_addr_off\[2\] _1630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Left_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3585__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4782__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5706_ _2059_ _2743_ _2745_ net843 _2748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6686_ _0259_ clknet_leaf_92_core_clock immu_1.high_addr_off\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3898_ _1391_ _1561_ _1562_ _1563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6594__CLK clknet_leaf_24_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_2501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_2512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5637_ _2708_ _0338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input370_I ic1_wb_adr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5568_ _2669_ _0308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input64_I c0_o_req_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold130 dmmu0.page_table\[13\]\[12\] net864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold141 dmmu1.page_table\[11\]\[1\] net875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4519_ _1852_ _2033_ _2035_ dmmu1.page_table\[14\]\[3\] _2039_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold152 dmmu1.page_table\[8\]\[5\] net886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5499_ _1976_ _2206_ _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold163 immu_0.page_table\[11\]\[3\] net897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold174 immu_1.page_table\[8\]\[8\] net908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold185 immu_1.page_table\[2\]\[3\] net919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold196 dmmu0.page_table\[6\]\[5\] net930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_10_980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4837__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Left_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7169_ net168 net624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6039__A1 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3273__A1 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3488__C _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6937__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3120__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4525__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4525__B2 dmmu1.page_table\[14\]\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_11__f_core_clock clknet_3_5_0_core_clock clknet_4_11__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6317__CLK clknet_leaf_70_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4289__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3187__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6467__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3264__A1 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4461__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4870_ _1812_ _2242_ _2244_ net767 _2251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5005__A2 _2336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3821_ immu_0.page_table\[4\]\[3\] immu_0.page_table\[5\]\[3\] immu_0.page_table\[6\]\[3\]
+ immu_0.page_table\[7\]\[3\] _1487_ _1455_ _1488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__4213__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3567__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6540_ _0113_ clknet_leaf_26_core_clock immu_0.page_table\[7\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3752_ _1308_ _1420_ _1421_ net663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_1293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_2068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6471_ _0044_ clknet_leaf_31_core_clock dmmu0.page_table\[8\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3683_ _1348_ net378 _1356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5422_ _2451_ _2582_ _2584_ net743 _2586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3319__A2 _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5353_ _2545_ _0217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4304_ _1907_ _0615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5284_ _2505_ _0188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3178__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4235_ net207 _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_78_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_2017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4166_ _1807_ _0577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_65_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3117_ _0866_ _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4097_ _1348_ net383 _1755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4047__A3 _1706_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5244__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input216_I dcache_mem_o_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3048_ _0824_ net474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6807_ _0380_ clknet_leaf_50_core_clock dmmu1.page_table\[11\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3809__S _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _1994_ _2316_ _2318_ net866 _2334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4755__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6738_ _0311_ clknet_leaf_46_core_clock dmmu1.page_table\[15\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6669_ _0242_ clknet_leaf_107_core_clock immu_0.high_addr_off\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_1407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4507__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5704__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5180__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3544__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output435_I net435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5483__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3494__A1 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output602_I net602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3246__A1 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4994__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3341__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4020_ net659 _1680_ _1681_ net672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_75_1636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5226__A2 _2469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3237__A1 _0982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5971_ _2849_ _2890_ _2892_ net1003 _2902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4922_ _2283_ _0048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_2078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3332__S1 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4853_ _1779_ _2205_ _2240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_7_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3804_ _1470_ _1471_ _1446_ _1472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4784_ _1812_ _2191_ _2193_ immu_0.page_table\[12\]\[6\] _2200_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6523_ _0096_ clknet_leaf_6_core_clock immu_0.page_table\[9\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3735_ _1404_ _1405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_42_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6454_ _0027_ clknet_leaf_38_core_clock dmmu0.page_table\[9\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3666_ _0814_ net320 _1326_ _1343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5405_ _2575_ _0239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5162__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6385_ _0767_ clknet_leaf_73_core_clock immu_1.page_table\[10\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6632__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3597_ net220 _1219_ _1299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_60_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input166_I c1_o_req_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5336_ _1977_ _2155_ _2535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_41_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6111__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5267_ _1811_ _2486_ _2488_ immu_0.page_table\[1\]\[6\] _2495_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_input333_I ic1_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4218_ _1850_ _0586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3476__A1 net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5198_ _2452_ _0155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input27_I c0_o_mem_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4149_ _1777_ _1792_ _1794_ immu_0.page_table\[11\]\[0\] _1795_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5217__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4425__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4976__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3323__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4728__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5925__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3400__A1 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5153__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3467__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4664__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3801__I _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3314__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6505__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5392__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5664__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6655__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3520_ net123 _1255_ _1257_ _1258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_68_1473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3451_ _1187_ _1190_ _1191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6170_ _3015_ _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3382_ net1 net53 _1119_ _1123_ _0841_ _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA_clkbuf_leaf_67_core_clock_I clknet_4_12__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1072 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5121_ _2405_ _0125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5052_ _2364_ _0097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_1381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4003_ _1633_ _1665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4407__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4958__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5954_ _2893_ _0470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4958__B2 dmmu0.page_table\[7\]\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4905_ _2273_ _2261_ _2263_ net768 _2274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5885_ _2047_ _2835_ _2837_ dmmu1.page_table\[8\]\[11\] _2853_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4836_ _2231_ _0014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5907__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4767_ _1972_ _2154_ _2189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3158__I _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input283_I ic0_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6506_ _0079_ clknet_leaf_7_core_clock immu_0.page_table\[10\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3718_ immu_0.page_table\[1\]\[0\] _1385_ _1387_ _1388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_44_997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4698_ _2065_ _2139_ _2142_ immu_1.page_table\[10\]\[5\] _2148_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_82_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5135__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6437_ _0010_ clknet_leaf_31_core_clock dmmu0.page_table\[10\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3649_ _0814_ net316 _1326_ _1330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5686__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_1844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6368_ _0750_ clknet_leaf_77_core_clock immu_1.page_table\[12\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5319_ _2461_ _2516_ _2518_ net1025 _2525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6299_ _0681_ clknet_leaf_85_core_clock immu_1.page_table\[1\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput305 ic0_mem_data[6] net305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3792__S1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3822__S _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold12 immu_0.page_table\[14\]\[7\] net746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput316 ic0_wb_adr[1] net316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput327 ic0_wb_sel[1] net327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5438__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold23 dmmu1.page_table\[10\]\[7\] net757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput338 ic1_mem_data[16] net338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput349 ic1_mem_data[26] net349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3449__A1 net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold34 dmmu0.page_table\[8\]\[5\] net768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold45 immu_1.page_table\[15\]\[5\] net779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4646__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold56 dmmu0.page_table\[6\]\[10\] net790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold67 dmmu1.page_table\[3\]\[7\] net801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4110__A2 net325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold78 immu_0.page_table\[8\]\[0\] net812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold89 dmmu1.page_table\[5\]\[1\] net823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_19_1604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6528__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_3_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5071__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5610__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3621__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6678__CLK clknet_leaf_40_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4177__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Left_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_1602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_9 net393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5126__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_2082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4627__I net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4101__A2 net380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5670_ _2682_ _2725_ _2727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_13_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4621_ net208 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_26_953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4552_ _2059_ _2053_ _2055_ immu_1.page_table\[15\]\[2\] _2060_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3471__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3503_ _0876_ _1240_ _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_23_core_clock clknet_4_4__leaf_core_clock clknet_leaf_23_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_13_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4483_ _1824_ _2014_ _2016_ immu_1.page_table\[3\]\[0\] _2017_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_1118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6222_ _0604_ clknet_leaf_86_core_clock immu_1.page_table\[7\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5668__A2 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3434_ dmmu0.page_table\[12\]\[10\] dmmu0.page_table\[13\]\[10\] dmmu0.page_table\[14\]\[10\]
+ dmmu0.page_table\[15\]\[10\] _0871_ _0866_ _1174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3679__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4876__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6153_ _1854_ _3000_ _3002_ immu_1.page_table\[8\]\[4\] _3007_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3774__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3365_ _0860_ _1107_ _0861_ _0821_ _1108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_5104_ _2394_ _0119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6084_ _2966_ _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3296_ dmmu1.page_table\[4\]\[5\] dmmu1.page_table\[5\]\[5\] dmmu1.page_table\[6\]\[5\]
+ dmmu1.page_table\[7\]\[5\] _0888_ _0901_ _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__6093__A2 _2957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5035_ _2265_ _2352_ _2354_ immu_0.page_table\[9\]\[1\] _2356_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input129_I c1_o_mem_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5840__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_2761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_85_2772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_2783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6820__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_2636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Left_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6986_ _0559_ clknet_leaf_79_core_clock immu_1.page_table\[8\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_81_2647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5937_ _2794_ _2873_ _2875_ net781 _2883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3603__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4800__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3089__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_2079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_62_core_clock clknet_4_14__leaf_core_clock clknet_leaf_62_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_5_1370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5868_ _2788_ _2836_ _2838_ net1034 _2843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input94_I c0_sr_bus_data_o[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5356__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4819_ _2220_ _0008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6970__CLK clknet_leaf_62_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3206__I1 _0953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3817__S _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5799_ _2803_ _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_66_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_2576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_2587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6200__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3214__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4331__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3552__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput102 c0_sr_bus_data_o[7] net102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput113 c1_o_instr_long_addr[3] net113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput124 c1_o_mem_addr[15] net124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6350__CLK clknet_leaf_63_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput135 c1_o_mem_data[10] net135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4619__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput146 c1_o_mem_data[6] net146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_51_1750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput157 c1_o_mem_high_addr[7] net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_51_1761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output515_I net515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput168 c1_o_req_addr[13] net168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4447__I net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput179 c1_o_req_addr[9] net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4095__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3842__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Right_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4182__I net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3070__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4910__I _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3453__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput609 net609 ic0_wb_i_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3526__I _1262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_28_Right_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_58_1948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_1959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3205__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4858__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3756__S1 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3150_ net121 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_20_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6075__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3081_ net162 net57 _0842_ _0843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6843__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Right_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6840_ _0413_ clknet_leaf_45_core_clock dmmu1.page_table\[9\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5035__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6993__CLK clknet_leaf_94_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6771_ _0344_ clknet_leaf_99_core_clock dmmu0.page_table\[5\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3983_ _1348_ _1645_ _1646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_1100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5188__I _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5722_ _2105_ _2742_ _2744_ dmmu1.page_table\[12\]\[10\] _2756_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5338__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5653_ _2717_ _0345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6223__CLK clknet_leaf_94_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _2091_ _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5889__A2 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Right_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5584_ _2677_ _0316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4535_ net199 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xhold301 immu_0.page_table\[6\]\[5\] net1035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4561__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold312 dmmu1.page_table\[7\]\[7\] net1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold323 dmmu1.page_table\[2\]\[1\] net1057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_2451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold334 immu_0.page_table\[4\]\[10\] net1068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold345 dmmu0.page_table\[14\]\[7\] net1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_70_2304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4466_ _2006_ _0678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6373__CLK clknet_leaf_96_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold356 dmmu1.page_table\[10\]\[9\] net1090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4849__B1 _2225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold367 dmmu0.page_table\[12\]\[11\] net1101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6205_ _0587_ clknet_leaf_96_core_clock immu_1.page_table\[9\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4313__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3417_ net154 dmmu1.long_off_reg\[4\] _1157_ _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_0_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3747__S1 _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7185_ net404 net657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4397_ _1852_ _1957_ _1959_ net859 _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input246_I dcache_wb_adr[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6136_ _1771_ _0809_ _0819_ _2995_ _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_77_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3348_ _0912_ _1088_ _1090_ _1091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_5_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6067_ net200 _2940_ _2942_ net828 _2956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4077__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Right_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3279_ _0882_ _1023_ _1024_ _0952_ _1025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_68_2244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_2709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5018_ _2345_ _0082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_68_2255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_2266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5577__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6969_ _0542_ clknet_leaf_60_core_clock dmmu1.page_table\[0\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_1380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_64_Right_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4001__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6716__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4552__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output632_I net632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3107__A3 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5501__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6866__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_73_Right_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6057__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4068__A1 net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5265__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5804__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3815__A1 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3130__I3 _0874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5017__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_82_Right_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4240__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5740__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3977__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput406 net406 c0_i_core_int_sreg[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_65_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput417 net417 c0_i_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4320_ _1918_ _0620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput428 net428 c0_i_req_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput439 net439 c0_i_req_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4251_ _1839_ _1873_ _1874_ _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_38_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3202_ _0864_ _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4182_ net104 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_38_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I c0_o_c_data_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3133_ _0860_ _0861_ _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_37_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3064_ net229 _0831_ _0833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_54_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6823_ _0396_ clknet_leaf_52_core_clock dmmu1.page_table\[10\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5559__A1 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6754_ _0327_ clknet_leaf_35_core_clock dmmu0.page_table\[6\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3966_ net7 immu_0.high_addr_off\[2\] _1629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_2_2052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5705_ _2747_ _0367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6739__CLK clknet_leaf_46_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_2085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6685_ _0258_ clknet_leaf_104_core_clock icache_arbiter.o_sel_sig vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4782__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3897_ _1385_ immu_0.page_table\[14\]\[5\] _1562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_76_2502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_2513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input196_I c1_sr_bus_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5636_ _1811_ _2699_ _2701_ dmmu0.page_table\[5\]\[6\] _2708_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_85_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_0__f_core_clock clknet_3_0_0_core_clock clknet_4_0__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_72_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5567_ _2059_ _2664_ _2666_ net950 _2669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_83_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6889__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold120 dmmu1.page_table\[10\]\[6\] net854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input363_I ic1_wb_adr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4518_ _2038_ _0698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold131 dmmu1.page_table\[13\]\[5\] net865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold142 dmmu1.page_table\[6\]\[9\] net876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_83_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold153 immu_0.page_table\[9\]\[10\] net887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5498_ _2628_ _0279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold164 dmmu1.page_table\[9\]\[5\] net898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input57_I c0_o_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold175 dmmu0.page_table\[4\]\[3\] net909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold186 dmmu1.page_table\[4\]\[6\] net920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4449_ _1995_ _0672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_1379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold197 immu_0.page_table\[7\]\[2\] net931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7168_ net167 net623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6039__A2 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6119_ _2847_ _2975_ _2977_ net821 _2986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7099_ net354 net507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_1718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5798__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_2105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6269__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4525__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5722__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_36_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4289__A1 _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5238__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__A1 _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3820_ _1369_ _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_24_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4213__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_1261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3751_ _1337_ net234 _1421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5961__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6470_ _0043_ clknet_leaf_31_core_clock dmmu0.page_table\[8\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3682_ _1353_ _1354_ _1355_ net682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_70_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5421_ _2585_ _0245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5352_ _2461_ _2536_ _2538_ net831 _2545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4303_ net209 _1894_ _1897_ immu_1.page_table\[0\]\[9\] _1907_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5283_ _1796_ _2502_ _2504_ immu_0.page_table\[0\]\[1\] _2505_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3714__I _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5477__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4234_ _1862_ _0590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6411__CLK clknet_leaf_112_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4165_ _1806_ _1792_ _1794_ net976 _1807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_65_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3116_ net16 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4096_ _1747_ _1753_ _1754_ net675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3047_ net221 _0822_ _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_78_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input111_I c1_o_instr_long_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input209_I c1_sr_bus_data_o[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6561__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6806_ _0379_ clknet_leaf_50_core_clock dmmu1.page_table\[11\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_74_core_clock_I clknet_4_11__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4998_ _2333_ _0074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_2095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_2114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3949_ _1611_ _1612_ net669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4755__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6737_ _0310_ clknet_leaf_46_core_clock dmmu1.page_table\[15\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_1968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6668_ _0241_ clknet_leaf_107_core_clock immu_0.high_addr_off\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5619_ _2697_ _0331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5704__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6599_ _0172_ clknet_leaf_17_core_clock immu_0.page_table\[2\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3825__S _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5180__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3560__S _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_2014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5640__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4994__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5943__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4190__I net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4054__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6434__CLK clknet_leaf_112_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4682__A1 _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6584__CLK clknet_leaf_24_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ _2901_ _0478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4921_ _1996_ _2260_ _2262_ dmmu0.page_table\[8\]\[12\] _2283_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4852_ _2239_ _0022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3803_ immu_1.page_table\[0\]\[2\] immu_1.page_table\[1\]\[2\] immu_1.page_table\[2\]\[2\]
+ immu_1.page_table\[3\]\[2\] _1435_ _1469_ _1471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4783_ _2199_ _0802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5196__I _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6522_ _0095_ clknet_leaf_7_core_clock immu_0.page_table\[9\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3734_ net366 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_42_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4033__C net705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6453_ _0026_ clknet_leaf_31_core_clock dmmu0.page_table\[9\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3665_ _1302_ net374 _1342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5404_ immu_0.high_addr_off\[2\] _1800_ _2572_ _2575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3548__I0 net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6384_ _0766_ clknet_leaf_97_core_clock immu_1.page_table\[10\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_1490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3596_ _1298_ net416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5335_ _2534_ _0210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input159_I c1_o_mem_req vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5266_ _2494_ _0181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6111__A1 _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6927__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4217_ _1849_ _1841_ _1843_ immu_1.page_table\[9\]\[2\] _1850_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_1794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5197_ _2451_ _2447_ _2449_ net841 _2452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5870__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input326_I ic0_wb_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4148_ _1793_ _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_39_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4079_ _1434_ _1738_ _1739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4425__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4976__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5925__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4728__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5153__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4664__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3303__B _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4185__I net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6169__A1 _2029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5392__A2 _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_13_core_clock clknet_4_3__leaf_core_clock clknet_leaf_13_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_0_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3450_ _1157_ _1188_ _1189_ _1190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3381_ net48 dmmu0.long_off_reg\[3\] _1122_ _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_21_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _2271_ _2398_ _2400_ immu_0.page_table\[6\]\[4\] _2405_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5051_ _2330_ _2352_ _2354_ net800 _2364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4002_ _1422_ _1663_ _1664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5852__B1 _2820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3213__B _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4407__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5604__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5953_ _2776_ _2890_ _2892_ dmmu1.page_table\[5\]\[0\] _2893_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4958__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4904_ _1808_ _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_52_core_clock clknet_4_13__leaf_core_clock clknet_leaf_52_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5884_ _2852_ _0441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4835_ _1806_ _2224_ _2226_ dmmu0.page_table\[10\]\[4\] _2231_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5907__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4766_ _2188_ _0796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3394__A1 net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4591__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6505_ _0078_ clknet_leaf_7_core_clock immu_0.page_table\[10\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3717_ _1386_ _1385_ _1387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4697_ _2147_ _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input276_I ic0_mem_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6436_ _0009_ clknet_leaf_108_core_clock immu_0.page_table\[13\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3648_ _1302_ net370 _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6183__I1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4343__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6367_ _0749_ clknet_leaf_63_core_clock immu_1.page_table\[12\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3579_ net226 _1204_ _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5318_ _2524_ _0203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6298_ _0680_ clknet_leaf_82_core_clock immu_1.page_table\[1\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput306 ic0_mem_data[7] net306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput317 ic0_wb_adr[2] net317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xhold13 immu_0.page_table\[8\]\[4\] net747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput328 ic0_wb_stb net328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5249_ _2483_ _0175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold24 dmmu0.page_table\[10\]\[9\] net758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput339 ic1_mem_data[17] net339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold35 immu_1.page_table\[6\]\[7\] net769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold46 dmmu0.page_table\[5\]\[5\] net780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4646__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold57 dmmu0.page_table\[5\]\[7\] net791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold68 dmmu1.page_table\[2\]\[6\] net802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold79 immu_1.page_table\[14\]\[7\] net813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_leaf_91_core_clock clknet_4_8__leaf_core_clock clknet_leaf_91_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5071__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5829__I _2820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3621__A2 net267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output495_I net495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5374__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output662_I net662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4009__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5126__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_2050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3084__I _0844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6087__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_13__f_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6622__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4620_ _2100_ _0738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3376__A1 _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4551_ _1848_ _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3502_ dmmu0.page_table\[8\]\[12\] dmmu0.page_table\[9\]\[12\] dmmu0.page_table\[10\]\[12\]
+ dmmu0.page_table\[11\]\[12\] _0863_ net16 _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3471__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4482_ _2015_ _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_41_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6221_ _0603_ clknet_leaf_87_core_clock immu_1.page_table\[7\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4325__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3433_ _1171_ _1172_ _0877_ _1173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5668__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4876__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3679__A2 net377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6152_ _3006_ _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3364_ net47 dmmu0.long_off_reg\[2\] _1106_ _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_TAPCELL_ROW_72_2390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5103_ _2330_ _2382_ _2384_ immu_0.page_table\[7\]\[9\] _2394_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_57_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6083_ _2790_ _2958_ _2960_ dmmu1.page_table\[1\]\[5\] _2966_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3295_ _1013_ _1040_ net524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__4628__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5034_ _2355_ _0088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_0_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_13_core_clock_I clknet_4_3__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5053__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6985_ _0558_ clknet_leaf_74_core_clock immu_1.page_table\[8\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_81_2637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_2648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5936_ _2882_ _0463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4800__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3603__A2 net382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5867_ _2842_ _0434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input393_I inner_wb_i_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5356__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4818_ _1819_ _2208_ _2210_ immu_0.page_table\[13\]\[9\] _2220_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5798_ _2682_ _2801_ _2803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input87_I c0_sr_bus_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4564__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4749_ _1800_ _2175_ _2177_ immu_0.page_table\[14\]\[2\] _2180_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6419_ _0801_ clknet_leaf_111_core_clock immu_0.page_table\[12\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3214__S1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput103 c0_sr_bus_data_o[8] net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_60_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput114 c1_o_instr_long_addr[4] net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput125 c1_o_mem_addr[1] net125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7104__I net389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput136 c1_o_mem_data[11] net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4619__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5816__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput147 c1_o_mem_data[7] net147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_51_1751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput158 c1_o_mem_long_mode net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_51_1762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput169 c1_o_req_addr[14] net169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4095__A2 net246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output508_I net508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6645__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1072 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6795__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3453__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_0_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3205__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4858__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3080_ _0841_ _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5283__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_4_core_clock_I clknet_4_1__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3982_ _1378_ _1639_ _1644_ _1382_ _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6770_ _0343_ clknet_leaf_42_core_clock dmmu0.page_table\[5\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3597__A1 net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_3_core_clock clknet_4_1__leaf_core_clock clknet_leaf_3_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_45_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5721_ _2755_ _0375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_1183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_79_core_clock_I clknet_4_11__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ dmmu0.long_off_reg\[0\] _1777_ _2716_ _2717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5338__A2 _2535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3349__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4603_ _1912_ _2089_ _2091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4546__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5889__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5583_ _2105_ _2663_ _2665_ dmmu1.page_table\[15\]\[10\] _2677_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4534_ _2046_ _0706_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold302 immu_1.page_table\[8\]\[6\] net1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6518__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_2430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold313 immu_0.page_table\[2\]\[9\] net1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold324 dmmu1.page_table\[5\]\[10\] net1058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold335 dmmu0.page_table\[5\]\[3\] net1069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_7_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4465_ _1854_ _1999_ _2001_ immu_1.page_table\[1\]\[4\] _2006_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xhold346 immu_1.page_table\[7\]\[1\] net1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold357 dmmu0.page_table\[1\]\[5\] net1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4849__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold368 dmmu1.page_table\[13\]\[6\] net1102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3416_ _1155_ _1127_ _1156_ _1157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6204_ _0586_ clknet_leaf_97_core_clock immu_1.page_table\[9\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7184_ net403 net656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4396_ _1962_ _0652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3521__A1 net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4548__I _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6135_ _2994_ mem_dcache_arb.select _2995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3347_ _0906_ _1089_ _1090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6668__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input141_I c1_o_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input239_I dcache_wb_adr[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6066_ _2955_ _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3278_ _0865_ dmmu0.page_table\[0\]\[4\] _1024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5017_ _2273_ _2337_ _2339_ immu_0.page_table\[10\]\[5\] _2345_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_68_2245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5577__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6968_ _0541_ clknet_leaf_58_core_clock dmmu1.page_table\[0\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5919_ _1873_ _1909_ _2031_ _2872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6899_ _0472_ clknet_leaf_54_core_clock dmmu1.page_table\[5\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_40_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6198__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output458_I net458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_53_1802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3107__A4 net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5501__A2 _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_81_core_clock_I clknet_4_10__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3512__A1 net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output625_I net625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5265__A1 _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3815__A2 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3371__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5017__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3311__B _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3123__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3579__A1 net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4776__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4240__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3537__I _1268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5740__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput407 net407 c0_i_core_int_sreg[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_50_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput418 net418 c0_i_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3751__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput429 net429 c0_i_req_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_65_1285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6810__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4250_ net188 net181 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3201_ _0930_ _0935_ _0947_ _0949_ net521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_38_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4700__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4181_ _1818_ _0581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3132_ _0864_ _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_38_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_2000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6960__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3063_ _0832_ net481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5199__I _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_2120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6822_ _0395_ clknet_leaf_49_core_clock dmmu1.page_table\[10\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5559__A2 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6753_ _0326_ clknet_leaf_34_core_clock dmmu0.page_table\[6\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3965_ net107 _1617_ _1627_ _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5704_ _2057_ _2743_ _2745_ net759 _2747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3896_ _1463_ immu_0.page_table\[15\]\[5\] _1561_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6684_ _0257_ clknet_leaf_101_core_clock dmmu0.page_table\[2\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6340__CLK clknet_leaf_73_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3990__A1 net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4519__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5635_ _2707_ _0337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_76_2503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input189_I c1_sr_bus_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5566_ _2668_ _0307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold110 immu_1.page_table\[13\]\[7\] net844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_2059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold121 dmmu1.page_table\[11\]\[10\] net855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4517_ _1849_ _2033_ _2035_ dmmu1.page_table\[14\]\[2\] _2038_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold132 dmmu0.page_table\[14\]\[11\] net866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5497_ net95 _2612_ _2614_ dmmu0.page_table\[4\]\[12\] _2628_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold143 immu_1.page_table\[4\]\[8\] net877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6490__CLK clknet_leaf_99_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold154 dmmu0.page_table\[10\]\[0\] net888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold165 immu_1.page_table\[7\]\[7\] net899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input356_I ic1_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold176 dmmu0.page_table\[6\]\[11\] net910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4448_ _1994_ _1978_ _1981_ dmmu0.page_table\[0\]\[11\] _1995_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold187 immu_1.page_table\[13\]\[1\] net921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5495__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold198 dmmu0.page_table\[10\]\[7\] net932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3182__I _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4379_ _1864_ _1942_ _1944_ net895 _1952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7167_ net166 net622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6039__A3 _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6118_ _2985_ _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7098_ net352 net505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6049_ _2786_ _2941_ _2943_ net1018 _2947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3558__S _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_1785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3981__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6833__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3733__A1 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4289__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6983__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5238__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3820__I _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3344__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4997__B1 _2318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4749__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4213__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3750_ _1401_ _1403_ _1419_ _1350_ _1420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_40_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5961__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3681_ _1337_ net253 _1355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5174__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5420_ _2444_ _2582_ _2584_ net1000 _2585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_40_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3724__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5351_ _2544_ _0216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4921__B1 _2262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4302_ _1906_ _0614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5282_ _2500_ _2502_ _2504_ _1386_ _0187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_43_2081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5477__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4233_ _1861_ _1841_ _1843_ net1109 _1862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4164_ _1805_ _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3115_ _0864_ _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4826__I _2225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4095_ _1535_ net246 _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4988__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3046_ _0823_ net467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6706__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input104_I c0_sr_bus_data_o[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6805_ _0378_ clknet_leaf_69_core_clock dmmu1.page_table\[12\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4997_ _2332_ _2316_ _2318_ dmmu0.page_table\[14\]\[10\] _2333_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6856__CLK clknet_leaf_100_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6736_ _0309_ clknet_leaf_48_core_clock dmmu1.page_table\[15\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_2058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3948_ _1306_ net240 _1612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3963__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6667_ _0240_ clknet_leaf_107_core_clock immu_0.high_addr_off\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3879_ _1440_ _1543_ _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5618_ net95 _2680_ _2683_ net809 _2697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4507__A3 _2029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5704__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6598_ _0171_ clknet_leaf_18_core_clock immu_0.page_table\[2\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5549_ _2527_ _2647_ _2649_ dmmu0.page_table\[3\]\[8\] _2658_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7112__I net403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6386__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5640__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4443__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4054__S1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6729__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4682__A2 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_2085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4920_ _2282_ _0047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_42_core_clock clknet_4_12__leaf_core_clock clknet_leaf_42_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_1734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_18_core_clock_I clknet_4_4__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4851_ _1996_ _2223_ _2225_ net806 _2239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4198__A1 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3802_ immu_1.page_table\[8\]\[2\] immu_1.page_table\[9\]\[2\] immu_1.page_table\[10\]\[2\]
+ immu_1.page_table\[11\]\[2\] _1435_ _1469_ _1470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_28_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4782_ _1809_ _2191_ _2193_ immu_0.page_table\[12\]\[5\] _2199_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_55_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3945__A1 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6521_ _0094_ clknet_leaf_6_core_clock immu_0.page_table\[9\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3733_ _0813_ _1402_ _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_67_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5147__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6452_ _0025_ clknet_leaf_17_core_clock dmmu0.page_table\[9\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3664_ _1339_ _1340_ _1341_ net678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5698__A1 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3548__I1 net31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _2574_ _0238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6259__CLK clknet_leaf_90_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3595_ net219 _1219_ _1298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6383_ _0765_ clknet_leaf_74_core_clock immu_1.page_table\[10\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_2007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5334_ _1996_ _2515_ _2517_ dmmu0.page_table\[12\]\[12\] _2534_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5265_ _1808_ _2486_ _2488_ immu_0.page_table\[1\]\[5\] _2494_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6111__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4122__A1 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4216_ _1848_ _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5196_ _1796_ _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5870__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_81_core_clock clknet_4_10__leaf_core_clock clknet_leaf_81_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4147_ _1771_ _1791_ _1793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input221_I dcache_mem_o_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3308__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input319_I ic0_wb_adr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4078_ immu_1.page_table\[12\]\[10\] immu_1.page_table\[13\]\[10\] immu_1.page_table\[14\]\[10\]
+ immu_1.page_table\[15\]\[10\] _1404_ _1540_ _1738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_74_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5622__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4425__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3029_ mem_dcache_arb.req1_pending net159 _0810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5386__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5925__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6719_ _0292_ clknet_leaf_11_core_clock dmmu0.page_table\[13\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_1176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7107__I net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_20_core_clock_I clknet_4_4__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4361__A1 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output440_I net440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput590 net590 ic0_mem_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__4113__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6167__B _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4664__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_9_core_clock_I clknet_4_1__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3927__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6401__CLK clknet_leaf_112_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3545__I _1272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3380_ _1106_ _1120_ _1121_ _1122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_20_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6551__CLK clknet_leaf_26_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5050_ _2363_ _0096_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4001_ _1502_ _1657_ _1662_ _1408_ _1663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__5852__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5604__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4407__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5455__I1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5952_ _2891_ _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_48_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4903_ _2272_ _0040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5883_ _2851_ _2835_ _2837_ dmmu1.page_table\[8\]\[10\] _2852_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4834_ _2230_ _0013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5907__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3918__A1 net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4765_ _1821_ _2174_ _2176_ net917 _2188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_2107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6504_ _0077_ clknet_leaf_3_core_clock immu_0.page_table\[10\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4591__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3716_ net737 _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4696_ _2063_ _2139_ _2142_ net840 _2147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6435_ _0008_ clknet_leaf_112_core_clock immu_0.page_table\[13\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3647_ _1325_ _1327_ _1328_ net660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input171_I c1_o_req_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4343__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input269_I dcache_wb_o_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6366_ _0748_ clknet_leaf_76_core_clock immu_1.page_table\[12\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3578_ _1289_ net422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5317_ _2459_ _2516_ _2518_ dmmu0.page_table\[12\]\[5\] _2524_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6297_ _0679_ clknet_leaf_82_core_clock immu_1.page_table\[1\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput307 ic0_mem_data[8] net307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput318 ic0_wb_adr[3] net318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xhold14 immu_0.page_table\[7\]\[8\] net748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput329 ic0_wb_we net329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5248_ _2332_ _2469_ _2471_ net998 _2483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold25 dmmu1.page_table\[12\]\[1\] net759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input32_I c0_o_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_86_core_clock_I clknet_4_10__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold36 dmmu1.page_table\[12\]\[11\] net770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4646__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold47 dmmu1.page_table\[6\]\[7\] net781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_58_1611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold58 dmmu1.page_table\[5\]\[7\] net792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold69 dmmu0.page_table\[6\]\[8\] net803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_58_1622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5179_ _2439_ _0149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5071__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6424__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3909__A1 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output488_I net488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4009__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_2046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4885__A2 _1972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1946 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_8__f_core_clock clknet_3_4_0_core_clock clknet_4_8__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_24_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_56_1888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6087__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5834__A1 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5598__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_1862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6011__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3984__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4573__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3376__A2 _1112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4550_ _2058_ _0710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_52_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3501_ _1237_ _1238_ _0875_ _1239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4481_ _1912_ _2013_ _2015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6220_ _0602_ clknet_leaf_86_core_clock immu_1.page_table\[7\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4325__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3759__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3432_ dmmu0.page_table\[0\]\[10\] dmmu0.page_table\[1\]\[10\] dmmu0.page_table\[2\]\[10\]
+ dmmu0.page_table\[3\]\[10\] _0871_ _0867_ _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_81_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4876__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3363_ _1077_ _1104_ _1105_ _1106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6151_ _1851_ _3000_ _3002_ net942 _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_72_2380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_2391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5102_ _2393_ _0118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3294_ net19 _1015_ _1016_ _1039_ _0884_ _1040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6082_ _2965_ _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_1519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5033_ _2258_ _2352_ _2354_ immu_0.page_table\[9\]\[0\] _2355_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3931__S0 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6984_ _0557_ clknet_leaf_81_core_clock immu_1.page_table\[8\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_85_2796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_2638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5935_ _2792_ _2873_ _2875_ net817 _2882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3064__A1 net229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4261__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4800__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5866_ _2786_ _2836_ _2838_ dmmu1.page_table\[8\]\[3\] _2842_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6597__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4817_ _2219_ _0007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5797_ _2801_ _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_1_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input386_I inner_ext_irq vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4564__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3367__A2 _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4748_ _2179_ _0787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3998__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_2589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4679_ _2135_ _0762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_1_Right_1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5513__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6418_ _0800_ clknet_leaf_109_core_clock immu_0.page_table\[12\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6349_ _0731_ clknet_leaf_62_core_clock immu_1.page_table\[13\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6069__A1 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4010__S _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput104 c0_sr_bus_data_o[9] net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput115 c1_o_instr_long_addr[5] net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput126 c1_o_mem_addr[2] net126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_42_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4619__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5816__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput137 c1_o_mem_data[12] net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_51_1741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput148 c1_o_mem_data[8] net148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_51_1752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput159 c1_o_mem_req net159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_51_1763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7120__I net59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3055__A1 net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_2050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4555__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4858__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5658__I1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5283__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3294__A1 net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4491__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3294__B2 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7030__I net386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5035__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3981_ _1378_ _1641_ _1643_ _1644_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4243__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5720_ _2103_ _2743_ _2745_ net811 _2755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_57_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3597__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5991__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5651_ _2715_ _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_2_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4602_ _2089_ _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4546__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3349__A2 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5582_ _2676_ _0315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4533_ _1870_ _2032_ _2034_ dmmu1.page_table\[14\]\[10\] _2046_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold303 immu_1.page_table\[11\]\[9\] net1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_74_2431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold314 dmmu0.page_table\[8\]\[10\] net1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_2442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold325 immu_0.page_table\[13\]\[3\] net1059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4464_ _2005_ _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold336 dmmu1.page_table\[5\]\[12\] net1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_68_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold347 immu_1.page_table\[14\]\[2\] net1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_68_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_2306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4849__A2 _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold358 immu_0.page_table\[5\]\[5\] net1092 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_68_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_2317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6203_ _0585_ clknet_leaf_81_core_clock immu_1.page_table\[9\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold369 immu_0.page_table\[8\]\[6\] net1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3415_ net153 dmmu1.long_off_reg\[3\] _1156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7183_ net402 net655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4395_ _1849_ _1957_ _1959_ net1066 _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_1242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6134_ mem_dcache_arb.transfer_active _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3521__A2 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3346_ dmmu1.page_table\[8\]\[7\] dmmu1.page_table\[9\]\[7\] dmmu1.page_table\[10\]\[7\]
+ dmmu1.page_table\[11\]\[7\] _0898_ _0909_ _1089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_42_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6065_ net199 _2940_ _2942_ net973 _2955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3277_ dmmu0.page_table\[1\]\[4\] _1023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input134_I c1_o_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5016_ _2344_ _0081_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_68_2246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3285__A1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input301_I ic0_mem_data[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6967_ _0540_ clknet_leaf_57_core_clock dmmu1.page_table\[0\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5918_ _2871_ _0456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6898_ _0471_ clknet_leaf_55_core_clock dmmu1.page_table\[5\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5849_ _2831_ _0427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5734__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_1803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7115__I net391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6612__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_1315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output520_I net520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5265__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4473__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3371__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5017__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_2101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4225__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_17_Left_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3123__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4776__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3579__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3200__A1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput408 net408 c0_i_irq vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput419 net419 c0_i_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3751__A2 net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_26_Left_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_1248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3553__I _1276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3200_ _0948_ _0862_ _0842_ _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4700__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4180_ _1817_ _1792_ _1794_ immu_0.page_table\[11\]\[8\] _1818_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3131_ _0862_ _0880_ _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3062_ net228 _0831_ _0832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_56_1901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3267__A1 net124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3267__B2 _1012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Left_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_2110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6821_ _0394_ clknet_leaf_49_core_clock dmmu1.page_table\[10\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_2121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5559__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4767__A1 _1972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6752_ _0325_ clknet_leaf_16_core_clock dmmu0.page_table\[6\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3964_ _0813_ _1626_ _1627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5703_ _2746_ _0366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6683_ _0256_ clknet_leaf_101_core_clock dmmu0.page_table\[2\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3895_ _1558_ _1559_ _1367_ _1560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4519__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5634_ _1808_ _2699_ _2701_ net780 _2707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4519__B2 dmmu1.page_table\[14\]\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5716__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_2504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5192__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5565_ _2057_ _2664_ _2666_ net860 _2668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6635__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Left_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold100 dmmu0.page_table\[3\]\[7\] net834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4516_ _2037_ _0697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold111 immu_0.page_table\[3\]\[9\] net845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold122 dmmu1.page_table\[12\]\[0\] net856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold133 dmmu0.page_table\[15\]\[4\] net867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5496_ _2627_ _0278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold144 immu_1.page_table\[7\]\[3\] net878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold155 dmmu1.page_table\[9\]\[1\] net889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4447_ net94 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xhold166 immu_0.page_table\[5\]\[6\] net900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold177 immu_0.page_table\[15\]\[10\] net911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input251_I dcache_wb_adr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold188 immu_0.page_table\[8\]\[3\] net922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_22_1613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5495__A2 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_25_core_clock_I clknet_4_5__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold199 dmmu0.page_table\[8\]\[2\] net933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input349_I ic1_mem_data[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7166_ net165 net621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6785__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4378_ _1951_ _0645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6117_ _1863_ _2975_ _2977_ net1042 _2985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3329_ dmmu0.page_table\[0\]\[6\] dmmu0.page_table\[1\]\[6\] dmmu0.page_table\[2\]\[6\]
+ dmmu0.page_table\[3\]\[6\] _0872_ _0941_ _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7097_ net351 net504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6048_ _2946_ _0511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3258__A1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3839__S _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5955__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4930__A1 _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4694__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5238__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4997__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3344__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_32_core_clock clknet_4_7__leaf_core_clock clknet_leaf_32_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4749__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6658__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3680_ _1350_ net323 _1326_ _1354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5174__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ _2459_ _2536_ _2538_ net871 _2544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4921__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4301_ net208 _1894_ _1897_ immu_1.page_table\[0\]\[8\] _1906_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5281_ _2503_ _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_49_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5477__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4232_ _1860_ _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_62_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3488__A1 _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_71_core_clock clknet_4_9__leaf_core_clock clknet_leaf_71_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4163_ net99 _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_39_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3114_ _0863_ _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4094_ _1750_ _1751_ _1752_ _1360_ _1753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__4437__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3232__B _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4988__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3045_ net214 _0822_ _0823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6804_ _0377_ clknet_leaf_43_core_clock dmmu1.page_table\[12\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5937__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4996_ net93 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_11_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6735_ _0308_ clknet_leaf_48_core_clock dmmu1.page_table\[15\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3947_ net659 _1594_ _1610_ _1611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3412__A1 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6666_ _0239_ clknet_leaf_109_core_clock immu_0.high_addr_off\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input299_I ic0_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3878_ immu_1.page_table\[8\]\[5\] immu_1.page_table\[9\]\[5\] immu_1.page_table\[10\]\[5\]
+ immu_1.page_table\[11\]\[5\] _1404_ _1540_ _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_60_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5617_ _2696_ _0330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6597_ _0170_ clknet_leaf_22_core_clock immu_0.page_table\[2\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5548_ _2657_ _0300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input62_I c0_o_req_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5479_ _2455_ _2613_ _2615_ net909 _2619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_6_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4676__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7149_ net404 net619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5640__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6800__CLK clknet_leaf_44_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3403__A1 _1119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_2011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6105__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5758__I _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4850_ _2238_ _0021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3801_ _1410_ _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_74_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4781_ _2198_ _0801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6520_ _0093_ clknet_leaf_4_core_clock immu_0.page_table\[9\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3732_ _1370_ _1382_ _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6451_ _0024_ clknet_leaf_30_core_clock dmmu0.page_table\[9\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5147__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3663_ _1337_ net249 _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5402_ immu_0.high_addr_off\[1\] _1797_ _2572_ _2574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5698__A2 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6382_ _0764_ clknet_leaf_79_core_clock immu_1.page_table\[10\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3594_ _1297_ net415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_1323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3227__B _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5333_ _2533_ _0209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5264_ _2493_ _0180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4215_ net202 _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4122__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5195_ _2450_ _0154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5870__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4146_ _1791_ _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3881__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3308__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6823__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4077_ _1440_ _1736_ _1737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input214_I dcache_mem_o_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5622__A2 _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3028_ mem_dcache_arb.req0_pending net54 _0809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3633__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3389__S _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5386__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6973__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4979_ _2322_ _0066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6718_ _0291_ clknet_leaf_14_core_clock dmmu0.page_table\[13\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6649_ _0222_ clknet_leaf_12_core_clock dmmu0.page_table\[15\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6203__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4361__A2 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6353__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput580 net580 dcache_wb_i_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput591 net591 ic0_mem_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_output433_I net433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7123__I net68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output600_I net600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_1145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3927__A2 _1590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_2052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5301__A1 net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3561__I _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6846__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4000_ _1415_ _1659_ _1661_ _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_79_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5852__A2 _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3863__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5604__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ _1770_ _2889_ _2891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3615__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6996__CLK clknet_leaf_97_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4812__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ _2271_ _2261_ _2263_ dmmu0.page_table\[8\]\[4\] _2272_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5882_ net198 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_47_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4833_ _1803_ _2224_ _2226_ net858 _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5368__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6226__CLK clknet_leaf_89_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4764_ _2187_ _0795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6503_ _0076_ clknet_leaf_10_core_clock dmmu0.page_table\[14\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3715_ _1384_ _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_55_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4591__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4695_ _2146_ _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6434_ _0007_ clknet_leaf_112_core_clock immu_0.page_table\[13\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3646_ _1306_ net231 _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_1950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4343__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6365_ _0747_ clknet_leaf_76_core_clock immu_1.page_table\[12\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3577_ net225 _1204_ _1289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input164_I c1_o_req_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5316_ _2523_ _0202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6296_ _0678_ clknet_leaf_83_core_clock immu_1.page_table\[1\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput308 ic0_mem_data[9] net308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5247_ _2482_ _0174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput319 ic0_wb_adr[4] net319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xhold15 immu_0.page_table\[4\]\[0\] net749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold26 immu_1.page_table\[6\]\[4\] net760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input331_I ic1_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold37 dmmu0.page_table\[6\]\[6\] net771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold48 dmmu0.page_table\[15\]\[3\] net782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold59 immu_1.page_table\[15\]\[9\] net793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5178_ _2275_ _2430_ _2432_ net966 _2439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input25_I c0_o_mem_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ _1775_ net658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_2010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3606__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3847__S _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4031__A1 _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6719__CLK clknet_leaf_11_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7118__I net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5531__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6869__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_2058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_1889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6087__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4098__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5295__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5834__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3845__A1 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5598__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6249__CLK clknet_leaf_90_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3757__S _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4940__I _2298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6011__A2 _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4022__A1 net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6399__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3456__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3500_ dmmu0.page_table\[4\]\[12\] dmmu0.page_table\[5\]\[12\] dmmu0.page_table\[6\]\[12\]
+ dmmu0.page_table\[7\]\[12\] _0863_ _0866_ _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_53_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4480_ _2013_ _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_40_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3208__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4325__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3431_ dmmu0.page_table\[4\]\[10\] dmmu0.page_table\[5\]\[10\] dmmu0.page_table\[6\]\[10\]
+ dmmu0.page_table\[7\]\[10\] _0871_ _0867_ _1171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3759__S1 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5771__I _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6150_ _3005_ _0554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3362_ net46 dmmu0.long_off_reg\[1\] _1105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_57_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_2370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _2328_ _2382_ _2384_ net748 _2393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_72_2392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6081_ _2788_ _2958_ _2960_ dmmu1.page_table\[1\]\[4\] _2965_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4089__A1 net116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3293_ _0879_ _1021_ _1026_ _1031_ _1038_ _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_20_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5032_ _2353_ _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3836__A1 _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3931__S1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5589__A1 _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6983_ _0556_ clknet_leaf_80_core_clock immu_1.page_table\[8\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_85_2786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5934_ _2881_ _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_66_2196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_2052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4261__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3064__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5865_ _2841_ _0433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4816_ _1817_ _2208_ _2210_ net1020 _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5796_ _1829_ _2031_ _2801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_69_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4747_ _1797_ _2175_ _2177_ net892 _2179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4564__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5761__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3998__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input281_I ic0_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input379_I ic1_wb_cyc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4678_ _2103_ _2123_ _2125_ net1037 _2135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6417_ _0799_ clknet_leaf_110_core_clock immu_0.page_table\[12\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5513__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3629_ _0812_ net271 _1318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_1600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6348_ _0730_ clknet_leaf_71_core_clock immu_1.page_table\[14\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1092 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6069__A2 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput105 c0_sr_bus_we net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6279_ _0661_ clknet_leaf_39_core_clock dmmu0.page_table\[0\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput116 c1_o_instr_long_addr[6] net116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput127 c1_o_mem_addr[3] net127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5816__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput138 c1_o_mem_data[13] net138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_51_1742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput149 c1_o_mem_data[9] net149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_51_1753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3827__A1 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3055__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_32_core_clock_I clknet_4_7__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5752__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6691__CLK clknet_4_8__leaf_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4307__A2 net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5591__I _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4491__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_1802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3980_ _1368_ _1642_ _1643_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4243__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5440__B1 _2583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5991__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4794__A2 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_2060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5650_ _1975_ _2570_ _2715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _1828_ _1839_ _2028_ _2089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_72_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4546__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5581_ _2103_ _2664_ _2666_ dmmu1.page_table\[15\]\[9\] _2676_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_1611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4532_ _2045_ _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold304 immu_0.page_table\[4\]\[2\] net1038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold315 immu_0.page_table\[2\]\[8\] net1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4463_ _1851_ _1999_ _2001_ immu_1.page_table\[1\]\[3\] _2005_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xhold326 dmmu1.page_table\[9\]\[12\] net1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_1920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold337 dmmu0.page_table\[14\]\[12\] net1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_46_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold348 dmmu1.page_table\[1\]\[3\] net1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_2307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6202_ _0584_ clknet_leaf_79_core_clock immu_1.page_table\[9\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3414_ net153 dmmu1.long_off_reg\[3\] _1155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
Xhold359 immu_1.page_table\[13\]\[8\] net1093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_42_1210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_2318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_15_Right_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_1953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7182_ net401 net654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_70_2329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4394_ _1961_ _0651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6133_ _1771_ _0810_ _0822_ _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_26_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3345_ _0896_ _1087_ _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5259__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6064_ _2954_ _0519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3276_ dmmu0.page_table\[2\]\[4\] dmmu0.page_table\[3\]\[4\] _0865_ _1022_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5015_ _2271_ _2337_ _2339_ immu_0.page_table\[10\]\[4\] _2344_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_2247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input127_I c1_o_mem_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6564__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_1648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_24_Right_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6966_ _0539_ clknet_leaf_59_core_clock dmmu1.page_table\[0\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5917_ _2049_ _2855_ _2857_ dmmu1.page_table\[7\]\[12\] _2871_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_33_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6897_ _0470_ clknet_leaf_55_core_clock dmmu1.page_table\[5\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _2529_ _2819_ _2821_ net1043 _2831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input92_I c0_sr_bus_data_o[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5734__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5779_ _2791_ _0397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_98_core_clock_I clknet_4_9__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_57_1940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3145__B _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_6__f_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6907__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output513_I net513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7131__I net61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4473__A1 net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_22_core_clock clknet_4_4__leaf_core_clock clknet_leaf_22_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_42_Right_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3028__A2 net54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4225__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5422__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4776__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3100__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_51_Right_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3200__A2 _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput409 net409 c0_i_mc_core_int vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6437__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5489__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4161__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4700__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_61_core_clock clknet_4_14__leaf_core_clock clknet_leaf_61_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_1596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3130_ _0869_ _0870_ _0873_ _0874_ _0877_ _0879_ _0880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_3061_ _0821_ _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7041__I net308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Right_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_2100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6820_ _0393_ clknet_leaf_50_core_clock dmmu1.page_table\[10\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_63_2111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6751_ _0324_ clknet_leaf_33_core_clock dmmu0.page_table\[6\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3963_ _1502_ _1620_ _1625_ _1408_ _1626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_46_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_2044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5702_ _2051_ _2743_ _2745_ net856 _2746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6682_ _0255_ clknet_leaf_100_core_clock dmmu0.page_table\[2\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3894_ immu_0.page_table\[0\]\[5\] immu_0.page_table\[1\]\[5\] immu_0.page_table\[2\]\[5\]
+ immu_0.page_table\[3\]\[5\] _1487_ _1390_ _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_85_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5633_ _2706_ _0336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4519__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5716__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5564_ _2667_ _0306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5192__A2 _2446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4515_ _1846_ _2033_ _2035_ dmmu1.page_table\[14\]\[1\] _2037_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold101 dmmu1.page_table\[1\]\[12\] net835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold112 dmmu0.page_table\[11\]\[11\] net846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold123 dmmu1.page_table\[1\]\[0\] net857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5495_ net94 _2612_ _2614_ dmmu0.page_table\[4\]\[11\] _2627_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold134 dmmu1.page_table\[10\]\[1\] net868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold145 dmmu1.page_table\[6\]\[11\] net879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold156 dmmu0.page_table\[11\]\[3\] net890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6141__A1 _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4446_ _1993_ _0671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold167 immu_0.page_table\[4\]\[8\] net901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_10_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold178 dmmu1.page_table\[6\]\[12\] net912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold189 dmmu1.page_table\[7\]\[3\] net923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7165_ net179 net635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4377_ _1861_ _1942_ _1944_ immu_1.page_table\[4\]\[6\] _1951_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_1625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input244_I dcache_wb_adr[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6116_ _2984_ _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3328_ dmmu0.page_table\[4\]\[6\] dmmu0.page_table\[5\]\[6\] dmmu0.page_table\[6\]\[6\]
+ dmmu0.page_table\[7\]\[6\] _0872_ _0941_ _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7096_ net350 net503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6047_ _2784_ _2941_ _2943_ dmmu1.page_table\[2\]\[2\] _2946_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3259_ dmmu1.page_table\[15\]\[4\] _1005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4455__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3412__C _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5400__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4207__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5955__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6949_ _0522_ clknet_leaf_58_core_clock dmmu1.page_table\[1\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3855__S _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3194__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4391__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7126__I net71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6132__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output630_I net630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4694__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4997__A2 _2316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4749__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5174__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3185__A1 net124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7036__I net303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4921__A2 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4300_ _1905_ _0613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5280_ _1895_ _2501_ _2503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6123__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4231_ net206 _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3488__A2 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4162_ _1804_ _0576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3113_ net15 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4093_ _1748_ _1731_ _1749_ _1752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4437__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5634__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3044_ _0821_ _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_56_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4988__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_1006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6803_ _0376_ clknet_leaf_69_core_clock dmmu1.page_table\[12\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5937__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3739__I net366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4995_ _2331_ _0073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6734_ _0307_ clknet_leaf_47_core_clock dmmu1.page_table\[15\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_2049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3946_ _1422_ _1605_ _1609_ _1610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_30_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3412__A2 _1147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6665_ _0238_ clknet_leaf_110_core_clock immu_0.high_addr_off\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3877_ _1434_ _1541_ _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_1359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input194_I c1_sr_bus_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5616_ net94 _2680_ _2683_ net910 _2696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_83_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6596_ _0169_ clknet_leaf_18_core_clock immu_0.page_table\[2\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4373__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6752__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5547_ _2463_ _2647_ _2649_ net834 _2657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input361_I ic1_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5478_ _2618_ _0269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input55_I c0_o_mem_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4429_ _1800_ _1979_ _1982_ dmmu0.page_table\[0\]\[2\] _1985_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3479__A2 _1214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4676__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7148_ net403 net618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7079_ net332 net485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_1810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6282__CLK clknet_leaf_40_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output678_I net678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3167__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6105__A1 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Left_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6625__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_2038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_16_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5919__A1 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3559__I _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_72_Left_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_1758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3800_ _1383_ _1460_ _1467_ _1468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_74_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4780_ _1806_ _2191_ _2193_ net1108 _2198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6775__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3731_ _1374_ _1379_ _1382_ _1400_ _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_28_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5774__I _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6450_ _0023_ clknet_leaf_31_core_clock dmmu0.page_table\[9\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3662_ _0814_ net319 _1326_ _1340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5147__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5401_ _2573_ _0237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4355__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6381_ _0763_ clknet_leaf_73_core_clock immu_1.page_table\[11\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5698__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3593_ net218 _1219_ _1297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_84_1482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ _1994_ _2515_ _2517_ net1101 _2533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_81_Left_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5263_ _1805_ _2486_ _2488_ immu_0.page_table\[1\]\[4\] _2493_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4658__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4214_ _1847_ _0585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5194_ _2444_ _2447_ _2449_ immu_0.page_table\[3\]\[0\] _2450_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4145_ _1781_ _1790_ _1791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_58_1827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4076_ immu_1.page_table\[8\]\[10\] immu_1.page_table\[9\]\[10\] immu_1.page_table\[10\]\[10\]
+ immu_1.page_table\[11\]\[10\] _1404_ _1540_ _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_78_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5083__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_2050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3633__A2 net258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input207_I c1_sr_bus_data_o[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5386__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4978_ _2267_ _2317_ _2319_ net832 _2322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3397__A1 net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6717_ _0290_ clknet_leaf_11_core_clock dmmu0.page_table\[13\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3929_ _1382_ _1587_ _1592_ _1593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA_clkbuf_leaf_37_core_clock_I clknet_4_7__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6648_ _0221_ clknet_leaf_11_core_clock dmmu0.page_table\[15\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6579_ _0152_ clknet_leaf_20_core_clock immu_0.page_table\[4\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4361__A3 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput570 net570 dcache_wb_i_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput581 net581 dcache_wb_i_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5846__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput592 net592 ic0_mem_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6648__CLK clknet_leaf_11_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_3_Left_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6798__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6023__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4585__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6177__I1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4888__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_2042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5950_ _2889_ _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4812__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3615__A2 net264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4901_ _1805_ _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_75_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ _2850_ _0440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4832_ _2229_ _0012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5368__A2 _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3379__A1 net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4763_ _1819_ _2175_ _2177_ immu_0.page_table\[14\]\[9\] _2187_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_83_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6502_ _0075_ clknet_leaf_12_core_clock dmmu0.page_table\[14\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3714_ _1369_ _1384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4694_ _2061_ _2139_ _2142_ net957 _2146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6433_ _0006_ clknet_leaf_111_core_clock immu_0.page_table\[13\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3645_ _0814_ net309 _1326_ _1327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3576_ _1288_ net421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6364_ _0746_ clknet_leaf_78_core_clock immu_1.page_table\[12\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5315_ _2457_ _2516_ _2518_ dmmu0.page_table\[12\]\[4\] _2523_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6295_ _0677_ clknet_leaf_90_core_clock immu_1.page_table\[1\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input157_I c1_o_mem_high_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput309 ic0_wb_adr[0] net309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_23_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5246_ _2330_ _2470_ _2472_ net1047 _2482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold16 immu_1.page_table\[12\]\[1\] net750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3303__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold27 immu_1.page_table\[11\]\[2\] net761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold38 dmmu0.page_table\[3\]\[9\] net772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5177_ _2438_ _0148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold49 immu_0.page_table\[9\]\[3\] net783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input324_I ic0_wb_adr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4128_ _0812_ net230 _1775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6940__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input18_I c0_o_mem_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4059_ immu_0.page_table\[8\]\[10\] immu_0.page_table\[9\]\[10\] immu_0.page_table\[10\]\[10\]
+ immu_0.page_table\[11\]\[10\] _1487_ _1390_ _1719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3606__A2 net328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3199__I _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4567__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4319__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5531__A2 _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7134__I net64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6470__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4098__A2 net329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5295__A1 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3845__A2 _1511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5047__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5598__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_2035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3153__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4558__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3456__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3081__I0 net162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3781__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3208__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3430_ _1170_ net530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6813__CLK clknet_leaf_44_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4730__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3361_ net46 dmmu0.long_off_reg\[1\] _1104_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_42_1425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7044__I net280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5100_ _2392_ _0117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6080_ _2964_ _0525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_72_2382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3292_ _0938_ _1034_ _1037_ _0878_ _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_72_2393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6963__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5031_ _2140_ _2351_ _2353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3392__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6982_ _0555_ clknet_leaf_74_core_clock immu_1.page_table\[8\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_85_2776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5933_ _2790_ _2873_ _2875_ net794 _2881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_66_2186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4261__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5864_ _2784_ _2836_ _2838_ net1039 _2841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6343__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4549__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4815_ _2218_ _0006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5795_ _2800_ _0404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4746_ _2178_ _0786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6493__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4677_ _2134_ _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_82_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input274_I dcache_wb_stb vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6416_ _0798_ clknet_leaf_1_core_clock immu_0.page_table\[12\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5513__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3628_ _1317_ net699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6347_ _0729_ clknet_leaf_78_core_clock immu_1.page_table\[14\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3559_ _1279_ net560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6069__A3 _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6278_ _0660_ clknet_leaf_95_core_clock immu_1.page_table\[6\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput106 c1_o_c_data_page net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput117 c1_o_instr_long_addr[7] net117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput128 c1_o_mem_addr[4] net128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput139 c1_o_mem_data[14] net139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5229_ _2473_ _0165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_51_1743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_1754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_12_core_clock clknet_4_3__leaf_core_clock clknet_leaf_12_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_1438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5202__I _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4788__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output493_I net493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7129__I net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6836__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3763__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4960__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6986__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3606__B net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_1160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_51_core_clock clknet_4_15__leaf_core_clock clknet_leaf_51_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_1789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_1808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6216__CLK clknet_leaf_91_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4491__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Left_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6366__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4243__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5440__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5991__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_2050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_2061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7039__I net306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4600_ _2088_ _0730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5580_ _2675_ _0314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_90_core_clock clknet_4_8__leaf_core_clock clknet_leaf_90_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_0_1260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ _1868_ _2033_ _2035_ dmmu1.page_table\[14\]\[9\] _2045_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_81_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold305 dmmu1.page_table\[8\]\[2\] net1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_83_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_2433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold316 immu_1.page_table\[4\]\[3\] net1050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4462_ _2004_ _0676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_74_2444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold327 immu_0.page_table\[5\]\[0\] net1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold338 dmmu0.page_table\[13\]\[0\] net1072 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6201_ _0583_ clknet_leaf_103_core_clock immu_0.page_table\[11\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3506__A1 net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold349 dmmu0.page_table\[7\]\[6\] net1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3413_ _1144_ _1153_ _0840_ _1154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_42_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_2319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4393_ _1846_ _1957_ _1959_ net1015 _1961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7181_ net400 net653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_1380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6132_ _1771_ _2992_ _2993_ _0548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_26_1987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3344_ dmmu1.page_table\[12\]\[7\] dmmu1.page_table\[13\]\[7\] dmmu1.page_table\[14\]\[7\]
+ dmmu1.page_table\[15\]\[7\] _0887_ _0909_ _1087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_61_1878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5259__A1 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3275_ _0948_ _1017_ _1020_ _0877_ _1021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6063_ _2851_ _2940_ _2942_ net1021 _2954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ _2343_ _0080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6709__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_1586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_2248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6965_ _0538_ clknet_leaf_53_core_clock dmmu1.page_table\[0\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6859__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5916_ _2870_ _0455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6896_ _0469_ clknet_leaf_68_core_clock dmmu1.page_table\[6\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_1384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5847_ _2830_ _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input391_I inner_wb_i_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5778_ _2790_ _2778_ _2780_ dmmu1.page_table\[10\]\[5\] _2791_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5734__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input85_I c0_sr_bus_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4729_ _2166_ _0781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3426__B net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6239__CLK clknet_leaf_82_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_1805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_1491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3356__S0 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6389__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4473__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5670__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output506_I net506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4225__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5422__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__A2 _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3984__A1 _1636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4933__B1 _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5489__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4161__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3060_ _0830_ net480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_1903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_2101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_2123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5777__I _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6750_ _0323_ clknet_leaf_33_core_clock dmmu0.page_table\[6\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3962_ _1415_ _1622_ _1624_ _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_58_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5701_ _2744_ _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_85_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6681_ _0254_ clknet_leaf_14_core_clock dmmu0.page_table\[2\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_1491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3893_ immu_0.page_table\[4\]\[5\] immu_0.page_table\[5\]\[5\] immu_0.page_table\[6\]\[5\]
+ immu_0.page_table\[7\]\[5\] _1487_ _1455_ _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_2_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5632_ _1805_ _2699_ _2701_ dmmu0.page_table\[5\]\[4\] _2706_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5716__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_2506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3727__A1 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5563_ _2051_ _2664_ _2666_ net913 _2667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_2007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4514_ _2036_ _0696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold102 dmmu1.page_table\[7\]\[9\] net836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold113 immu_0.page_table\[7\]\[0\] net847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5494_ _2626_ _0277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold124 dmmu0.page_table\[10\]\[3\] net858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold135 immu_1.page_table\[15\]\[0\] net869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4445_ _1821_ _1978_ _1981_ dmmu0.page_table\[0\]\[10\] _1993_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold146 immu_1.page_table\[10\]\[0\] net880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold157 dmmu1.page_table\[7\]\[0\] net891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6141__A2 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold168 dmmu1.page_table\[0\]\[1\] net902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_22_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold179 dmmu1.page_table\[15\]\[0\] net913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_10_952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7164_ net178 net634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4376_ _1950_ _0644_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6115_ _1860_ _2975_ _2977_ net929 _2984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3327_ _0934_ _1068_ _1070_ _1051_ _0841_ _1071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7095_ net349 net502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input237_I dcache_wb_adr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5101__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6046_ _2945_ _0510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3258_ _0931_ _1000_ _1003_ _0897_ _1004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_20_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3189_ _0877_ _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6681__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input404_I inner_wb_i_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6948_ _0521_ clknet_leaf_64_core_clock dmmu1.page_table\[2\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5955__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3966__A1 net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6879_ _0452_ clknet_leaf_61_core_clock dmmu1.page_table\[7\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5168__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4915__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4391__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4930__A3 _2286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4143__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5340__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_2_core_clock clknet_4_1__leaf_core_clock clknet_leaf_2_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_60_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4694__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5891__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output623_I net623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_109_core_clock clknet_4_0__leaf_core_clock clknet_leaf_109_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_40_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7142__I net397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3329__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_44_core_clock_I clknet_4_12__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6404__CLK clknet_leaf_110_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3709__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6554__CLK clknet_leaf_23_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6123__A2 _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4134__A1 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4230_ _1859_ _0589_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4161_ _1803_ _1792_ _1794_ net897 _1804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7052__I net289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3112_ _0860_ _0861_ _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4092_ _0813_ net107 _1751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5634__A1 _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4437__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3043_ _0819_ _0820_ _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_65_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_19_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6802_ _0375_ clknet_leaf_43_core_clock dmmu1.page_table\[12\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4994_ _2330_ _2317_ _2319_ dmmu0.page_table\[14\]\[9\] _2331_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5937__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3948__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6733_ _0306_ clknet_leaf_47_core_clock dmmu1.page_table\[15\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3945_ net107 _1608_ _1609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6664_ _0237_ clknet_leaf_109_core_clock immu_0.high_addr_off\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3876_ immu_1.page_table\[12\]\[5\] immu_1.page_table\[13\]\[5\] immu_1.page_table\[14\]\[5\]
+ immu_1.page_table\[15\]\[5\] _1404_ _1540_ _1541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_27_882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5615_ _2695_ _0329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3755__I _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6595_ _0168_ clknet_leaf_24_core_clock immu_0.page_table\[2\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4373__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input187_I c1_sr_bus_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5546_ _2656_ _0299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5477_ _2453_ _2613_ _2615_ net994 _2618_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input354_I ic1_mem_data[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4428_ _1984_ _0662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_6_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input48_I c0_o_mem_high_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4676__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7147_ net402 net617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4359_ _1870_ _1926_ _1928_ immu_1.page_table\[5\]\[10\] _1940_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7078_ net362 net515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_1508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_2018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6029_ _2847_ _2924_ _2926_ net999 _2935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4027__S _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3939__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6577__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_1859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5400__I1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6105__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5313__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5864__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_0_0_core_clock clknet_0_core_clock clknet_3_0_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5616__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_2011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5467__I1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_2017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_2077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_16_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5919__A2 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6041__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3776__S _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3730_ _1383_ _1393_ _1399_ _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_51_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_2050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3661_ _1302_ net373 _1339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7047__I net283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5400_ immu_0.high_addr_off\[0\] _1777_ _2572_ _2573_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4355__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3789__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6380_ _0762_ clknet_leaf_81_core_clock immu_1.page_table\[11\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3592_ _1296_ net414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5331_ _2532_ _0208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4107__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5262_ _2492_ _0179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4213_ _1846_ _1841_ _1843_ net1044 _1847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5193_ _2448_ _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_78_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4144_ _1789_ _1790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_23_1798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4075_ _1733_ _1734_ _1439_ _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5083__A2 _2381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4291__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_2095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input102_I c0_sr_bus_data_o[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4977_ _2321_ _0065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6716_ _0289_ clknet_leaf_14_core_clock dmmu0.page_table\[13\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3397__A2 net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3928_ _1378_ _1589_ _1591_ _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_46_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1946 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6647_ _0220_ clknet_leaf_15_core_clock dmmu0.page_table\[15\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3859_ _1368_ _1524_ _1525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_15_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5543__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6578_ _0151_ clknet_leaf_24_core_clock immu_0.page_table\[4\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5529_ _1976_ _2445_ _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_48_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5406__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6099__A1 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput560 net560 dcache_mem_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput571 net571 dcache_wb_i_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5846__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput582 net582 ic0_mem_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput593 net593 ic0_mem_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5205__I _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6023__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_2072 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4585__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4337__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4888__A2 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5065__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3076__A1 net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6742__CLK clknet_leaf_42_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4273__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4812__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4900_ _2270_ _0039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5880_ _2849_ _2836_ _2838_ dmmu1.page_table\[8\]\[9\] _2850_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4831_ _1800_ _2224_ _2226_ dmmu0.page_table\[10\]\[2\] _2229_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4762_ _2186_ _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6501_ _0074_ clknet_leaf_11_core_clock dmmu0.page_table\[14\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3713_ _1377_ _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_44_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4693_ _2145_ _0766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6432_ _0005_ clknet_leaf_0_core_clock immu_0.page_table\[13\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3644_ _1304_ _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5525__B1 _2631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6363_ _0745_ clknet_leaf_72_core_clock immu_1.page_table\[12\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3575_ net224 _1204_ _1288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_64_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5314_ _2522_ _0201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6294_ _0676_ clknet_leaf_90_core_clock immu_1.page_table\[1\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5828__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6272__CLK clknet_leaf_85_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5245_ _2481_ _0173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold17 immu_0.page_table\[11\]\[1\] net751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold28 immu_0.page_table\[14\]\[6\] net762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold39 immu_0.page_table\[10\]\[7\] net773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5176_ _2273_ _2430_ _2432_ immu_0.page_table\[4\]\[5\] _2438_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4127_ net659 _0816_ net565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_39_1024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_2012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input317_I ic0_wb_adr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4058_ _1383_ _1715_ _1717_ _1718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_75_1972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6005__A1 net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4567__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4319__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_41_core_clock clknet_4_6__leaf_core_clock clknet_leaf_41_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_1938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3164__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output536_I net536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5295__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6765__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7150__I net390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5047__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4255__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3153__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_2110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4558__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_80_core_clock clknet_4_10__leaf_core_clock clknet_leaf_80_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5507__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6295__CLK clknet_leaf_90_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4730__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3360_ _1096_ _1098_ _1100_ _1102_ _1103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_2372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3291_ _0882_ _1035_ _1036_ _0948_ _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA_clkbuf_4_1__f_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5030_ _2351_ _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3297__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3392__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3049__A1 net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3521__C _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6981_ _0554_ clknet_leaf_96_core_clock immu_1.page_table\[8\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_85_2766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5932_ _2880_ _0461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_85_2799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_2187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5863_ _2840_ _0432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4814_ _1815_ _2208_ _2210_ immu_0.page_table\[13\]\[7\] _2218_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4549__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5746__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5794_ _2049_ _2777_ _2779_ dmmu1.page_table\[10\]\[12\] _2800_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4745_ _1777_ _2175_ _2177_ net842 _2178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_56_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6638__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4676_ _2101_ _2123_ _2125_ net863 _2134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_1337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6415_ _0797_ clknet_leaf_109_core_clock immu_0.page_table\[12\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3627_ _1308_ net270 _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input267_I dcache_wb_o_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6346_ _0728_ clknet_leaf_76_core_clock immu_1.page_table\[14\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3558_ net160 net55 _0841_ _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6788__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6277_ _0659_ clknet_leaf_86_core_clock immu_1.page_table\[6\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3489_ net50 dmmu0.long_off_reg\[5\] _1228_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput107 c1_o_c_instr_long net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_55_1880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput118 c1_o_mem_addr[0] net118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5228_ _2444_ _2470_ _2472_ immu_0.page_table\[2\]\[0\] _2473_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3288__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput129 c1_o_mem_addr[5] net129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input30_I c0_o_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4485__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5159_ _2332_ _2413_ _2415_ net893 _2427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_32_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5029__A2 _2240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_49_core_clock_I clknet_4_13__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_32_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4237__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4788__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5985__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_1684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3460__A1 net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output486_I net486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3212__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3874__S _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4960__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3673__I _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7145__I net400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3279__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_101_core_clock_I clknet_4_2__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_1804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5440__A2 _2581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_2040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_2051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_2062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_core_clock_I clknet_4_15__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4530_ _2044_ _0704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_1050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4461_ _1848_ _1999_ _2001_ immu_1.page_table\[1\]\[2\] _2004_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6153__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold306 immu_1.page_table\[13\]\[0\] net1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold317 dmmu1.page_table\[3\]\[1\] net1051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7055__I net292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold328 dmmu1.page_table\[8\]\[6\] net1062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold339 immu_1.page_table\[8\]\[2\] net1073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6200_ _0582_ clknet_leaf_5_core_clock immu_0.page_table\[11\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_1802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3412_ _0878_ _1147_ _1152_ _0883_ _1153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_7180_ net399 net652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_2309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4392_ _1960_ _0650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6131_ net559 _2991_ mem_dcache_arb.select _2993_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3343_ _1084_ _1085_ _0896_ _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_1999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5259__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6062_ _2953_ _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3274_ _0882_ _1018_ _1019_ _0952_ _1020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4467__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5013_ _2269_ _2337_ _2339_ net822 _2343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_68_2249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__CLK clknet_leaf_85_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3690__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_1797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_5_Right_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5967__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6964_ _0537_ clknet_leaf_58_core_clock dmmu1.page_table\[0\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3817__I0 net236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _2047_ _2855_ _2857_ dmmu1.page_table\[7\]\[11\] _2870_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3442__A1 net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6895_ _0468_ clknet_leaf_66_core_clock dmmu1.page_table\[6\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5846_ _2527_ _2819_ _2821_ dmmu0.page_table\[1\]\[8\] _2830_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5777_ _1857_ _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_20_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input384_I inner_disable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4728_ _1812_ _2157_ _2159_ immu_0.page_table\[15\]\[6\] _2166_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4942__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input78_I c0_sr_bus_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4659_ _2124_ _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_57_1920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_2035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6329_ _0711_ clknet_leaf_72_core_clock immu_1.page_table\[15\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5414__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3356__S1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_5_0_core_clock clknet_0_core_clock clknet_3_5_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5670__A2 _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3681__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6803__CLK clknet_leaf_69_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5422__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5186__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6953__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4933__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4933__B2 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5489__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4161__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6333__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5110__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6483__CLK clknet_leaf_32_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3961_ _1440_ _1623_ _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5700_ _2682_ _2742_ _2744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_70_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6680_ _0253_ clknet_leaf_40_core_clock dmmu0.page_table\[2\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3892_ net2 _1556_ _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_14_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5631_ _2705_ _0335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_1380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5562_ _2665_ _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_54_883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4513_ _1824_ _2033_ _2035_ dmmu1.page_table\[14\]\[0\] _2036_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold103 dmmu1.page_table\[11\]\[0\] net837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5493_ _2531_ _2612_ _2614_ dmmu0.page_table\[4\]\[10\] _2626_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold114 dmmu0.page_table\[12\]\[3\] net848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold125 immu_1.page_table\[6\]\[3\] net859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4444_ _1992_ _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold136 dmmu1.page_table\[15\]\[4\] net870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold147 dmmu0.page_table\[2\]\[9\] net881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold158 immu_0.page_table\[14\]\[1\] net892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4688__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6141__A3 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold169 dmmu1.page_table\[4\]\[3\] net903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7163_ net177 net633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4375_ _1858_ _1942_ _1944_ net948 _1950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3360__B1 _1100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6114_ _2983_ _0540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3326_ net151 dmmu1.long_off_reg\[1\] _1069_ _1070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7094_ net348 net501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6045_ _2782_ _2941_ _2943_ net1057 _2945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5101__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3257_ _0889_ _1001_ _1002_ _0902_ _1003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__6826__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input132_I c1_o_mem_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3188_ dmmu0.page_table\[8\]\[1\] dmmu0.page_table\[9\]\[1\] dmmu0.page_table\[10\]\[1\]
+ dmmu0.page_table\[11\]\[1\] _0872_ _0868_ _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3663__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4860__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6976__CLK clknet_leaf_105_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4093__B _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3415__A1 net153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _0520_ clknet_leaf_65_core_clock dmmu1.page_table\[2\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_27_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6878_ _0451_ clknet_leaf_57_core_clock dmmu1.page_table\[7\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5168__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _2820_ _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6206__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4915__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3718__A2 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6117__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4391__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5208__I _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6356__CLK clknet_leaf_63_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5340__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output449_I net449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3329__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3654__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__B1 _2225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3900__B _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4134__A2 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6849__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4160_ _1802_ _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_4_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_69_2300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3111_ net1 net53 _0861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4091_ _1748_ _1731_ _1749_ _1750_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_21_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5095__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5634__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3042_ mem_dcache_arb.select net559 _0820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput290 ic0_mem_data[21] net290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3645__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_19_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6801_ _0374_ clknet_leaf_45_core_clock dmmu1.page_table\[12\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4993_ net104 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6229__CLK clknet_leaf_82_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3101__I _0853_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3944_ net112 immu_1.high_addr_off\[2\] _1607_ _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__3948__A2 net240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6732_ _0305_ clknet_leaf_97_core_clock dmmu0.page_table\[3\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6663_ _0236_ clknet_leaf_102_core_clock dmmu0.page_table\[11\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3875_ _1410_ _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_74_989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5614_ _2531_ _2680_ _2683_ net790 _2695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6379__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6594_ _0167_ clknet_leaf_24_core_clock immu_0.page_table\[2\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4373__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5545_ _2461_ _2647_ _2649_ net851 _2656_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5476_ _2617_ _0268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4427_ _1797_ _1979_ _1982_ dmmu0.page_table\[0\]\[1\] _1984_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3771__I _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input347_I ic1_mem_data[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7146_ net401 net616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4358_ _1939_ _0637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3309_ _0938_ _1053_ _1054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7077_ net361 net514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4289_ _1848_ _1894_ _1897_ immu_1.page_table\[0\]\[2\] _1900_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6028_ _2934_ _0503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_1981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4833__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_1987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5561__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_2069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5313__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7153__I net393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5864__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5077__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5616__A2 _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3627__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_2007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5919__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6041__A2 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3486__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6521__CLK clknet_leaf_6_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3660_ _1335_ _1336_ _1338_ net677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3238__S0 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5001__B1 _2318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4355__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3591_ net217 _1219_ _1296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3789__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6671__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5330_ _2531_ _2515_ _2517_ net1002 _2532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_84_1495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3805__B _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4107__A2 net273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5261_ _1802_ _2486_ _2488_ immu_0.page_table\[1\]\[3\] _2492_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4212_ _1845_ _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5192_ _1980_ _2446_ _2448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4143_ _1769_ _1785_ _1788_ _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_4
X_4074_ immu_1.page_table\[0\]\[10\] immu_1.page_table\[1\]\[10\] immu_1.page_table\[2\]\[10\]
+ immu_1.page_table\[3\]\[10\] _1435_ _1469_ _1734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4291__A1 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4976_ _2265_ _2317_ _2319_ dmmu0.page_table\[14\]\[1\] _2321_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5240__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6715_ _0288_ clknet_leaf_28_core_clock dmmu0.page_table\[13\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_1114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3927_ _1368_ _1590_ _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3766__I _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input297_I ic0_mem_data[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6646_ _0219_ clknet_leaf_28_core_clock dmmu0.page_table\[15\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3858_ immu_0.page_table\[0\]\[4\] immu_0.page_table\[1\]\[4\] immu_0.page_table\[2\]\[4\]
+ immu_0.page_table\[3\]\[4\] _1463_ _1391_ _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_85_1226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3229__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5543__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3789_ immu_0.page_table\[8\]\[2\] immu_0.page_table\[9\]\[2\] immu_0.page_table\[10\]\[2\]
+ immu_0.page_table\[11\]\[2\] _1424_ _1455_ _1457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6577_ _0150_ clknet_leaf_22_core_clock immu_0.page_table\[4\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5528_ _2645_ _0292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_31_core_clock clknet_4_7__leaf_core_clock clknet_leaf_31_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input60_I c0_o_req_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6099__A2 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5459_ immu_1.high_addr_off\[3\] _1852_ _2603_ _2607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput550 net550 dcache_mem_i_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput561 net561 dcache_mem_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput572 net572 dcache_wb_i_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5846__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput583 net583 ic0_mem_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3857__A1 _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput594 net594 ic0_mem_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3857__B2 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7129_ net74 net597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5059__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_106_core_clock_I clknet_4_2__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4806__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6544__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6023__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4034__A1 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3468__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output683_I net683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_70_core_clock clknet_4_9__leaf_core_clock clknet_leaf_70_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7148__I net403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_56_core_clock_I clknet_4_14__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3076__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4273__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_83_2694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4830_ _2228_ _0011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4761_ _1817_ _2175_ _2177_ immu_0.page_table\[14\]\[8\] _2186_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_51_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3712_ _1381_ _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_43_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6500_ _0073_ clknet_leaf_15_core_clock dmmu0.page_table\[14\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4692_ _2059_ _2139_ _2142_ immu_1.page_table\[10\]\[2\] _2145_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_4_5__f_core_clock clknet_3_2_0_core_clock clknet_4_5__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_1508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3643_ _1302_ net363 _1325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6431_ _0004_ clknet_leaf_0_core_clock immu_0.page_table\[13\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5525__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6362_ _0744_ clknet_leaf_76_core_clock immu_1.page_table\[12\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3574_ _1287_ net420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5313_ _2455_ _2516_ _2518_ net848 _2522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6417__CLK clknet_leaf_110_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6293_ _0675_ clknet_leaf_82_core_clock immu_1.page_table\[1\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5289__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5828__A2 _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5244_ _2328_ _2470_ _2472_ net1049 _2481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold18 dmmu0.page_table\[13\]\[11\] net752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold29 immu_0.page_table\[9\]\[2\] net763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5175_ _2437_ _0147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_1615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4126_ net659 _0815_ net564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_58_1626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6567__CLK clknet_leaf_26_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _1368_ _1716_ _1717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input212_I dcache_mem_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6005__A2 _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4016__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4567__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4959_ _2310_ _0058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4319__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6629_ _0202_ clknet_leaf_33_core_clock dmmu0.page_table\[12\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_2011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output431_I net431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3550__I0 net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3180__B _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4255__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_2059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4558__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5507__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3355__B _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4730__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3290_ _0882_ dmmu0.page_table\[12\]\[4\] _1036_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_72_2373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_2384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3297__A2 _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Left_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3049__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6980_ _0553_ clknet_leaf_81_core_clock immu_1.page_table\[8\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4246__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5931_ _2788_ _2873_ _2875_ dmmu1.page_table\[6\]\[4\] _2880_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_2188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5862_ _2782_ _2836_ _2838_ net1014 _2840_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4813_ _2217_ _0005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4549__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5746__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5793_ _2799_ _0403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_84_870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4744_ _2176_ _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_16_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_78_Left_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4675_ _2133_ _0760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3626_ _1316_ net698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6414_ _0796_ clknet_leaf_108_core_clock immu_0.page_table\[14\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3265__B _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3557_ _1278_ net549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6345_ _0727_ clknet_leaf_63_core_clock immu_1.page_table\[14\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_1062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input162_I c1_o_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6276_ _0658_ clknet_leaf_87_core_clock immu_1.page_table\[6\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3488_ _0875_ _1224_ _1226_ _0878_ _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_55_1870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput108 c1_o_c_instr_page net108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5227_ _2471_ _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_55_1881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput119 c1_o_mem_addr[10] net119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_1734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4485__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5682__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5158_ _2426_ _0141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input23_I c0_o_mem_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4109_ _1535_ net255 _1764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4237__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5089_ _2267_ _2382_ _2384_ net931 _2387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5434__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5985__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4788__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_1696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4115__I _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3212__A2 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4960__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output479_I net479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6732__CLK clknet_leaf_97_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4173__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7161__I net175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6882__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3523__I0 _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_2041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5728__A1 _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_2063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6262__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_2560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_2571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ _2003_ _0675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_2424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6153__A1 _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold307 dmmu0.page_table\[5\]\[10\] net1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_46_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_2435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold318 dmmu1.page_table\[13\]\[2\] net1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold329 immu_1.page_table\[12\]\[6\] net1063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3411_ _1149_ _1151_ _0878_ _1152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_68_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4391_ _1824_ _1957_ _1959_ immu_1.page_table\[6\]\[0\] _1960_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6130_ net559 _0818_ _2991_ _2992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_0_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3342_ dmmu1.page_table\[4\]\[7\] dmmu1.page_table\[5\]\[7\] dmmu1.page_table\[6\]\[7\]
+ dmmu1.page_table\[7\]\[7\] _0898_ _0909_ _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_42_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6061_ _2849_ _2941_ _2943_ dmmu1.page_table\[2\]\[9\] _2953_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3273_ _0865_ dmmu0.page_table\[4\]\[4\] _1019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4467__A1 _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4011__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5012_ _2342_ _0079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_1732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3690__A2 net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6963_ _0536_ clknet_leaf_56_core_clock dmmu1.page_table\[0\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5967__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5914_ _2869_ _0454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6894_ _0467_ clknet_leaf_67_core_clock dmmu1.page_table\[6\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5845_ _2829_ _0425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4078__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5776_ _2789_ _0396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_40_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6755__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4727_ _2165_ _0780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4942__A2 _2298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input377_I ic1_wb_adr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4658_ _1912_ _2122_ _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_1146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput90 c0_sr_bus_addr[8] net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_1921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3609_ _1303_ _1305_ _1307_ net703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_57_1932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4589_ _2065_ _2075_ _2077_ net799 _2083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_3_7_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6328_ _0710_ clknet_leaf_76_core_clock immu_1.page_table\[15\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_1807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6259_ _0641_ clknet_leaf_90_core_clock immu_1.page_table\[4\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3681__A2 net253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6285__CLK clknet_leaf_41_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4630__A1 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Right_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output596_I net596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5186__A2 _2429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4933__A2 _2285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7156__I net164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Right_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5110__A2 _2397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6628__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5949__A1 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_2103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3960_ immu_1.page_table\[8\]\[7\] immu_1.page_table\[9\]\[7\] immu_1.page_table\[10\]\[7\]
+ immu_1.page_table\[11\]\[7\] _1441_ _1442_ _1623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_9_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6778__CLK clknet_leaf_104_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1072 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3891_ _1553_ _1554_ _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6171__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5630_ _1802_ _2699_ _2701_ net1069 _2705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_14_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_2101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3807__S0 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4924__A2 _2222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5561_ _2300_ _2663_ _2665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7066__I net406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4512_ _2034_ _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5492_ _2625_ _0276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold104 dmmu1.page_table\[1\]\[7\] net838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold115 immu_1.page_table\[15\]\[8\] net849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold126 dmmu1.page_table\[15\]\[1\] net860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4443_ _1819_ _1979_ _1982_ net754 _1992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_1600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold137 dmmu0.page_table\[15\]\[5\] net871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4688__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold148 dmmu0.page_table\[0\]\[5\] net882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold159 immu_0.page_table\[5\]\[10\] net893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4374_ _1949_ _0643_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7162_ net176 net632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_81_1092 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3325_ net150 dmmu1.long_off_reg\[0\] _1069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6113_ _1857_ _2975_ _2977_ net1013 _2983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7093_ net347 net500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6044_ _2944_ _0509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3256_ _0899_ dmmu1.page_table\[8\]\[4\] _1002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_2075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5101__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3112__A1 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3187_ dmmu0.page_table\[12\]\[1\] dmmu0.page_table\[13\]\[1\] dmmu0.page_table\[14\]\[1\]
+ dmmu0.page_table\[15\]\[1\] _0872_ _0868_ _0936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4860__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3663__A2 net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input125_I c1_o_mem_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6946_ _0519_ clknet_leaf_65_core_clock dmmu1.page_table\[2\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6877_ _0450_ clknet_leaf_56_core_clock dmmu1.page_table\[7\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5168__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5828_ _2682_ _2818_ _2820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input90_I c0_sr_bus_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3179__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4915__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5759_ _2031_ _2137_ _2777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_17_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6117__A1 _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5340__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3351__A1 net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold1_I ic0_wb_cyc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5628__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output511_I net511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3654__A2 net247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4851__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6920__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6053__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4603__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5800__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4367__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6300__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6450__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3110_ net53 _0859_ _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XTAP_TAPCELL_ROW_69_2301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4090_ net117 immu_1.high_addr_off\[7\] _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5095__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3041_ net559 _0818_ _0819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4973__I _2318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3645__A2 net309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput280 ic0_mem_data[12] net280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput291 ic0_mem_data[22] net291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_63_core_clock_I clknet_4_11__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6800_ _0373_ clknet_leaf_44_core_clock dmmu1.page_table\[12\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4992_ _2329_ _0072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_19_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6731_ _0304_ clknet_leaf_100_core_clock dmmu0.page_table\[3\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3943_ _1606_ _1549_ _1607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6662_ _0235_ clknet_leaf_12_core_clock dmmu0.page_table\[11\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3874_ _1537_ _1538_ _1416_ _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _2694_ _0328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6593_ _0166_ clknet_leaf_19_core_clock immu_0.page_table\[2\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3257__C _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5544_ _2655_ _0298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_21_core_clock clknet_4_4__leaf_core_clock clknet_leaf_21_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_5_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3581__A1 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5475_ _2451_ _2613_ _2615_ dmmu0.page_table\[4\]\[1\] _2617_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_83_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4426_ _1983_ _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3333__A1 net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7145_ net400 net615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4357_ _1868_ _1927_ _1929_ immu_1.page_table\[5\]\[9\] _1939_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input242_I dcache_wb_adr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3308_ dmmu0.page_table\[12\]\[5\] dmmu0.page_table\[13\]\[5\] dmmu0.page_table\[14\]\[5\]
+ dmmu0.page_table\[15\]\[5\] _0872_ _0868_ _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_7076_ net360 net513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4288_ _1899_ _0607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3239_ dmmu1.page_table\[8\]\[3\] dmmu1.page_table\[9\]\[3\] dmmu1.page_table\[10\]\[3\]
+ dmmu1.page_table\[11\]\[3\] _0889_ _0931_ _0986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6027_ _2794_ _2924_ _2926_ net801 _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_1802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4833__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4597__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6929_ _0502_ clknet_leaf_58_core_clock dmmu1.page_table\[3\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_60_core_clock clknet_4_14__leaf_core_clock clknet_leaf_60_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6323__CLK clknet_leaf_70_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4349__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5561__A2 _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Left_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output559_I net559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6473__CLK clknet_leaf_101_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5313__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4521__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5077__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3911__B _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3627__A2 net270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Left_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_1421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_16_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3202__I _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3486__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5001__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3238__S1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_41_Left_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6816__CLK clknet_leaf_69_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3590_ _1295_ net413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3563__A1 _1154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5260_ _2491_ _0178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3315__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6966__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4211_ net201 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_27_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5191_ _2446_ _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4142_ net105 _1786_ _1787_ _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XPHY_EDGE_ROW_50_Left_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4073_ immu_1.page_table\[4\]\[10\] immu_1.page_table\[5\]\[10\] immu_1.page_table\[6\]\[10\]
+ immu_1.page_table\[7\]\[10\] _1435_ _1469_ _1733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3174__S0 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4291__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6346__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4579__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4975_ _2320_ _0064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5240__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6714_ _0287_ clknet_leaf_33_core_clock dmmu0.page_table\[13\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3926_ immu_0.page_table\[8\]\[6\] immu_0.page_table\[9\]\[6\] immu_0.page_table\[10\]\[6\]
+ immu_0.page_table\[11\]\[6\] _1424_ _1371_ _1590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_73_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6645_ _0218_ clknet_leaf_33_core_clock dmmu0.page_table\[15\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3857_ _1408_ _1521_ _1522_ net107 _1301_ _1523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_27_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6496__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3229__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input192_I c1_sr_bus_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5543__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6576_ _0149_ clknet_leaf_22_core_clock immu_0.page_table\[4\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3788_ immu_0.page_table\[0\]\[2\] immu_0.page_table\[1\]\[2\] immu_0.page_table\[2\]\[2\]
+ immu_0.page_table\[3\]\[2\] _1424_ _1455_ _1456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_14_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4751__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5527_ net95 _2629_ _2631_ net864 _2645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6099__A3 _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput540 net540 dcache_mem_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5458_ _2606_ _0261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input53_I c0_o_mem_long_mode vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput551 net551 dcache_mem_i_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3306__A1 net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput562 net562 dcache_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput573 net573 dcache_wb_i_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4409_ _1868_ _1957_ _1959_ immu_1.page_table\[6\]\[9\] _1969_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput584 net584 ic0_mem_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_80_1894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput595 net595 ic0_mem_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5389_ _2565_ _0233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3857__A2 _1521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7128_ net73 net596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5059__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3731__B _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7059_ net296 net447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5502__I _2631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4806__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4034__A2 _1694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3468__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6839__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3093__I0 net129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6989__CLK clknet_leaf_73_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3906__B _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7164__I net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6219__CLK clknet_leaf_90_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6369__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4273__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_2695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4760_ _2185_ _0793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3711_ net385 _1380_ net2 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__3784__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4691_ _2144_ _0765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_1282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _0003_ clknet_leaf_111_core_clock immu_0.page_table\[13\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3642_ _1324_ net691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5525__A2 _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6361_ _0743_ clknet_leaf_63_core_clock immu_1.page_table\[12\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3573_ net223 _1204_ _1287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7074__I net358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_49_Right_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5312_ _2521_ _0200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6292_ _0674_ clknet_leaf_83_core_clock immu_1.page_table\[1\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5289__A1 _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5243_ _2480_ _0172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_1531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold19 immu_0.page_table\[8\]\[2\] net753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5174_ _2271_ _2430_ _2432_ net915 _2437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4125_ _1774_ net483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4056_ immu_0.page_table\[0\]\[10\] immu_0.page_table\[1\]\[10\] immu_0.page_table\[2\]\[10\]
+ immu_0.page_table\[3\]\[10\] _1370_ _1391_ _1716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_75_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_58_Right_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input205_I c1_sr_bus_data_o[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3777__I _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4016__A2 _1672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4958_ _2277_ _2299_ _2302_ dmmu0.page_table\[7\]\[7\] _2310_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1092 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3775__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3909_ _1377_ _1573_ _1574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_69_1734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4889_ _2262_ _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_69_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6628_ _0201_ clknet_leaf_29_core_clock dmmu0.page_table\[12\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_1789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_67_Right_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4724__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6559_ _0132_ clknet_leaf_7_core_clock immu_0.page_table\[5\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_2078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6511__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3550__I1 net32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Right_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_1738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4255__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7159__I net173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3310__S0 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_85_Right_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5507__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4191__A1 net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_2374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5930_ _2879_ _0460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_85_2779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_2189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5861_ _2839_ _0431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4812_ _1812_ _2208_ _2210_ net1086 _2217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5792_ _2047_ _2777_ _2779_ dmmu1.page_table\[10\]\[11\] _2799_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5746__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4954__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4743_ _2140_ _2174_ _2176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4674_ _2069_ _2123_ _2125_ net874 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3509__A1 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6413_ _0795_ clknet_leaf_0_core_clock immu_0.page_table\[14\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4706__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3625_ _1308_ net269 _1316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_24_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6344_ _0726_ clknet_leaf_76_core_clock immu_1.page_table\[14\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3556_ net140 net35 _0841_ _1278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6534__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6275_ _0657_ clknet_leaf_86_core_clock immu_1.page_table\[6\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3487_ _0877_ _1225_ _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_45_1096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_1860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input155_I c1_o_mem_high_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3368__S0 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput109 c1_o_icache_flush net109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5226_ _1980_ _2469_ _2471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_55_1882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4485__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5682__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6684__CLK clknet_leaf_101_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5157_ _2330_ _2414_ _2416_ net850 _2426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input322_I ic0_wb_adr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4108_ _1761_ _1762_ _1763_ net702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_32_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5088_ _2386_ _0111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5434__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input16_I c0_o_mem_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4237__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4039_ net10 immu_0.high_addr_off\[5\] _1699_ _1700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__3501__S _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5985__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3748__A1 _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4131__I _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4173__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5370__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3920__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5122__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_68_core_clock_I clknet_4_12__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3210__I net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5728__A2 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_2550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3366__B _1108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_2561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6153__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_2425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold308 dmmu1.page_table\[0\]\[7\] net1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold319 immu_1.page_table\[3\]\[4\] net1053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3410_ _0877_ _1150_ _1151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3211__I0 _0956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ _1958_ _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_46_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3341_ dmmu1.page_table\[0\]\[7\] dmmu1.page_table\[1\]\[7\] dmmu1.page_table\[2\]\[7\]
+ dmmu1.page_table\[3\]\[7\] _0898_ _0901_ _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3813__C _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6060_ _2952_ _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3272_ dmmu0.page_table\[5\]\[4\] _1018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_20_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I c0_o_instr_long_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4011__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5011_ _2267_ _2337_ _2339_ immu_0.page_table\[10\]\[2\] _2342_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_84_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_2011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6962_ _0535_ clknet_leaf_58_core_clock dmmu1.page_table\[0\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5967__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_2006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3978__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5913_ _2851_ _2855_ _2857_ dmmu1.page_table\[7\]\[10\] _2869_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6893_ _0466_ clknet_leaf_59_core_clock dmmu1.page_table\[6\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4216__I _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5844_ _1814_ _2819_ _2821_ dmmu0.page_table\[1\]\[7\] _2829_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4078__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4927__B1 _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5775_ _2788_ _2778_ _2780_ dmmu1.page_table\[10\]\[4\] _2789_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_20_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4726_ _1809_ _2157_ _2159_ immu_0.page_table\[15\]\[5\] _2165_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4657_ _2122_ _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_70_core_clock_I clknet_4_9__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input272_I dcache_wb_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3608_ _1306_ net274 _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput80 c0_sr_bus_addr[13] net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5352__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput91 c0_sr_bus_addr[9] net91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_1933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4588_ _2082_ _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3902__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6327_ _0709_ clknet_leaf_63_core_clock immu_1.page_table\[15\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_2059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3539_ _1269_ net555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3723__C _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6258_ _0640_ clknet_leaf_86_core_clock immu_1.page_table\[4\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ _2459_ _2447_ _2449_ immu_0.page_table\[3\]\[5\] _2460_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6189_ _1796_ _3026_ _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3969__A1 net8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3513__S0 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4630__A2 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output491_I net491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3186__B _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7172__I net109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3406__S _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5646__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_2006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_2240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5949__A2 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3504__S0 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3890_ _1553_ _1554_ _1555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_15_1658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3875__I _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3807__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4385__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5560_ _2663_ _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_83_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_2509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_11_core_clock clknet_4_3__leaf_core_clock clknet_leaf_11_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4511_ _1980_ _2032_ _2034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_79_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5491_ _2529_ _2613_ _2615_ dmmu0.page_table\[4\]\[9\] _2625_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold105 dmmu1.page_table\[6\]\[0\] net839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_78_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold116 immu_0.page_table\[5\]\[9\] net850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4442_ _1991_ _0669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold127 dmmu0.page_table\[15\]\[12\] net861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_10_900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold138 dmmu1.page_table\[14\]\[12\] net872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold149 dmmu1.page_table\[13\]\[0\] net883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4688__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5885__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7161_ net175 net631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4373_ _1855_ _1942_ _1944_ net1033 _1949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7082__I net335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6112_ _2982_ _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3324_ _1064_ _1065_ _1066_ _1067_ _0906_ _0912_ _1068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_7092_ net346 net499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6043_ _2776_ _2941_ _2943_ dmmu1.page_table\[2\]\[0\] _2944_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3255_ dmmu1.page_table\[9\]\[4\] _1001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__3115__I _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3743__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3186_ _0931_ _0934_ _0884_ _0935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4860__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input118_I c1_o_mem_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _0518_ clknet_leaf_60_core_clock dmmu1.page_table\[2\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6722__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_50_core_clock clknet_4_13__leaf_core_clock clknet_leaf_50_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5660__I1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _0449_ clknet_leaf_57_core_clock dmmu1.page_table\[7\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_27_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5827_ _2818_ _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_48_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5412__I1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3179__A2 _0927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6872__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ _1823_ _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5573__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input83_I c0_sr_bus_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4709_ _2153_ _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6117__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5689_ _2737_ _0361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4128__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3226__S _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3351__A2 net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5628__A1 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6252__CLK clknet_leaf_89_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output504_I net504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4851__A2 _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6053__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5800__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4367__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_2302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5095__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3040_ mem_dcache_arb.req1_pending net159 _0809_ _0817_ _0818_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_21_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6745__CLK clknet_leaf_69_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput270 dcache_wb_o_dat[8] net270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput281 ic0_mem_data[13] net281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput292 ic0_mem_data[23] net292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4991_ _2328_ _2317_ _2319_ dmmu0.page_table\[14\]\[8\] _2329_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_19_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6730_ _0303_ clknet_leaf_98_core_clock dmmu0.page_table\[3\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3942_ net111 immu_1.high_addr_off\[1\] _1606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6895__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6661_ _0234_ clknet_leaf_102_core_clock dmmu0.page_table\[11\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3873_ immu_1.page_table\[4\]\[5\] immu_1.page_table\[5\]\[5\] immu_1.page_table\[6\]\[5\]
+ immu_1.page_table\[7\]\[5\] _1435_ _1469_ _1538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_6_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7077__I net361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5612_ _2529_ _2681_ _2684_ net766 _2694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6592_ _0165_ clknet_leaf_20_core_clock immu_0.page_table\[2\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5543_ _2459_ _2647_ _2649_ net755 _2655_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_83_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5307__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3581__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5474_ _2616_ _0267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput700 net700 inner_wb_o_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5858__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4425_ _1777_ _1979_ _1982_ dmmu0.page_table\[0\]\[0\] _1983_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6275__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7144_ net399 net614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4356_ _1938_ _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3307_ _0934_ _1049_ _1050_ _1051_ _0841_ _1052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7075_ net359 net512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4287_ _1845_ _1894_ _1897_ immu_1.page_table\[0\]\[1\] _1899_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_input235_I dcache_wb_adr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6026_ _2933_ _0502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3238_ dmmu1.page_table\[12\]\[3\] dmmu1.page_table\[13\]\[3\] dmmu1.page_table\[14\]\[3\]
+ dmmu1.page_table\[15\]\[3\] _0889_ _0931_ _0985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_20_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4833__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3169_ _0907_ _0918_ _0919_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input402_I inner_wb_i_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6035__A1 net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4597__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6928_ _0501_ clknet_leaf_58_core_clock dmmu1.page_table\[3\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6859_ _0432_ clknet_leaf_50_core_clock dmmu1.page_table\[8\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4349__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6618__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output454_I net454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4521__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3955__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4521__B2 dmmu1.page_table\[14\]\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6768__CLK clknet_leaf_41_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output621_I net621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3911__C _1575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3260__A1 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5537__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5001__A2 _2316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_2097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6298__CLK clknet_leaf_82_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3563__A2 _1186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4210_ _1844_ _0584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3166__I2 dmmu1.page_table\[14\]\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _1789_ _2445_ _2446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_62_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4141_ net89 net88 net87 _1787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__6177__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4072_ net107 _1730_ _1731_ _1732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_78_1268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3174__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6017__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4974_ _2258_ _2317_ _2319_ dmmu0.page_table\[14\]\[0\] _2320_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_1_core_clock clknet_4_0__leaf_core_clock clknet_leaf_1_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5240__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3925_ _1375_ _1588_ _1589_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6713_ _0286_ clknet_leaf_16_core_clock dmmu0.page_table\[13\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3251__A1 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_108_core_clock clknet_4_0__leaf_core_clock clknet_leaf_108_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_50_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4224__I _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6644_ _0217_ clknet_leaf_16_core_clock dmmu0.page_table\[15\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3856_ net110 immu_1.high_addr_off\[0\] _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6575_ _0148_ clknet_leaf_27_core_clock immu_0.page_table\[4\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3787_ net313 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_67_1662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4751__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input185_I c1_sr_bus_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5526_ _2644_ _0291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6910__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5457_ immu_1.high_addr_off\[2\] _1849_ _2603_ _2606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput530 net530 dcache_mem_addr[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput541 net541 dcache_mem_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput552 net552 dcache_mem_i_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input352_I ic1_mem_data[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput563 net563 dcache_rst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4408_ _1968_ _0658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4503__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput574 net574 dcache_wb_i_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5388_ _2529_ _2553_ _2555_ net1005 _2565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput585 net585 ic0_mem_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input46_I c0_o_mem_high_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput596 net596 ic0_mem_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_7127_ net72 net595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4339_ _1824_ _1927_ _1929_ immu_1.page_table\[5\]\[0\] _1930_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5059__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7058_ net295 net446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4267__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4806__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6009_ _1874_ _1891_ _2030_ _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_69_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3242__A1 _0974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3093__I1 net24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6440__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6590__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_2046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7180__I net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_14__f_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3710_ net3 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3784__A2 _1427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4690_ _2057_ _2139_ _2142_ immu_1.page_table\[10\]\[1\] _2144_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_0_core_clock_I clknet_4_0__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3641_ _0812_ net262 _1324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6933__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6360_ _0742_ clknet_leaf_63_core_clock immu_1.page_table\[12\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3572_ _1286_ net419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5311_ _2453_ _2516_ _2518_ net1076 _2521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_3_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6291_ _0673_ clknet_leaf_101_core_clock dmmu0.page_table\[0\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_75_core_clock_I clknet_4_11__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5289__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5242_ _2463_ _2470_ _2472_ immu_0.page_table\[2\]\[7\] _2480_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3919__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4497__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5173_ _2436_ _0146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4124_ net213 _0831_ _1774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6313__CLK clknet_leaf_94_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 c0_o_c_data_page net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_78_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4055_ _1375_ _1714_ _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3847__I0 net237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5997__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_2097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3472__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6463__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input100_I c0_sr_bus_data_o[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4957_ _2309_ _0057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3908_ _1563_ _1566_ _1569_ _1572_ _1573_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3775__A2 _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4972__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4888_ _1980_ _2260_ _2262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_12_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4889__I _2262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6627_ _0200_ clknet_leaf_33_core_clock dmmu0.page_table\[12\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3839_ immu_1.page_table\[12\]\[3\] immu_1.page_table\[13\]\[3\] _1474_ _1506_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_2002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4724__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6558_ _0131_ clknet_leaf_9_core_clock immu_0.page_table\[6\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5509_ _2455_ _2630_ _2632_ net960 _2636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6489_ _0062_ clknet_leaf_13_core_clock dmmu0.page_table\[7\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6806__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_2017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4660__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3310__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7175__I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6336__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ _2776_ _2836_ _2838_ net941 _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4811_ _2216_ _0004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5791_ _2798_ _0402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4403__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4954__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4742_ _2174_ _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_31_1867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4673_ _2132_ _0759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_1919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6412_ _0794_ clknet_leaf_112_core_clock immu_0.page_table\[14\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3624_ _1315_ net697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4706__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5903__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6343_ _0725_ clknet_leaf_76_core_clock immu_1.page_table\[14\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3555_ _1277_ net548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3118__I _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6274_ _0656_ clknet_leaf_89_core_clock immu_1.page_table\[6\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3486_ dmmu0.page_table\[0\]\[11\] dmmu0.page_table\[1\]\[11\] dmmu0.page_table\[2\]\[11\]
+ dmmu0.page_table\[3\]\[11\] _0871_ _0866_ _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5225_ _2469_ _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_55_1861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3368__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_1883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6829__CLK clknet_leaf_69_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input148_I c1_o_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5682__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5156_ _2425_ _0140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_1758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3693__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4890__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4107_ _1535_ net273 _1763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5087_ _2265_ _2382_ _2384_ immu_0.page_table\[7\]\[1\] _2386_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_32_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5434__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input315_I ic0_wb_adr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4038_ _1666_ _1697_ _1698_ _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6979__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4642__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5989_ _2786_ _2907_ _2909_ net903 _2913_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6209__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3748__A2 _1417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6147__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5370__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4173__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3920__A2 _1583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5122__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3684__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3698__I _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_2043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5728__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_78_2551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_2090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_2573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_2426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold309 dmmu0.page_table\[1\]\[9\] net1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_2448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3340_ net152 dmmu1.long_off_reg\[2\] _1082_ _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_81_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3271_ dmmu0.page_table\[6\]\[4\] dmmu0.page_table\[7\]\[4\] _0872_ _1017_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5010_ _2341_ _0078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4872__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6185__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6961_ _0534_ clknet_leaf_64_core_clock dmmu1.page_table\[1\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3427__A1 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5912_ _2868_ _0453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_40_core_clock clknet_4_6__leaf_core_clock clknet_leaf_40_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6892_ _0465_ clknet_leaf_61_core_clock dmmu1.page_table\[6\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ _2828_ _0424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4927__A1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4927__B2 _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_1551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5774_ _1854_ _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_12_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6501__CLK clknet_leaf_11_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4725_ _2164_ _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4232__I _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4656_ _1826_ _1839_ _1874_ _2122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_82_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput70 c0_o_req_addr[5] net70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3607_ inner_wb_arbiter.o_sel_sig _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput81 c0_sr_bus_addr[14] net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5352__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ _2063_ _2075_ _2077_ immu_1.page_table\[14\]\[4\] _2082_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_57_1923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput92 c0_sr_bus_data_o[0] net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6651__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input265_I dcache_wb_o_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3538_ net146 net41 _1267_ _1269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6326_ _0708_ clknet_leaf_70_core_clock dmmu1.page_table\[14\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3292__B _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6257_ _0639_ clknet_leaf_84_core_clock immu_1.page_table\[4\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_10_Left_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3469_ _0907_ _1207_ _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5208_ _1808_ _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6188_ _1781_ _1788_ _2284_ _3026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_23_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3666__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5139_ _2258_ _2414_ _2416_ net1061 _2417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3418__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4615__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3513__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4630__A3 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output484_I net484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5646__A2 _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3657__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3930__B _1593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_2230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5949__A3 _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6071__A2 _2957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3504__S1 net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4082__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6524__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_2084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4510_ _2032_ _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_53_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6674__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ _2624_ _0275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_14_core_clock_I clknet_4_6__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold106 immu_1.page_table\[10\]\[4\] net840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5334__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4441_ _1817_ _1979_ _1982_ dmmu0.page_table\[0\]\[8\] _1991_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold117 dmmu0.page_table\[3\]\[6\] net851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_9_Right_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold128 dmmu1.page_table\[12\]\[7\] net862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold139 immu_1.page_table\[6\]\[8\] net873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7160_ net174 net630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4372_ _1948_ _0642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3896__A1 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6111_ _1854_ _2975_ _2977_ dmmu1.page_table\[0\]\[4\] _2982_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3323_ dmmu1.page_table\[8\]\[6\] dmmu1.page_table\[9\]\[6\] dmmu1.page_table\[10\]\[6\]
+ dmmu1.page_table\[11\]\[6\] _0888_ _0901_ _1067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_10_956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7091_ net345 net498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4001__B _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6042_ _2942_ _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3254_ dmmu1.page_table\[10\]\[4\] dmmu1.page_table\[11\]\[4\] _0908_ _1000_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3648__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4936__B _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4845__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3743__S1 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3185_ net124 _0932_ _0892_ _0933_ _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
XANTENNA__4227__I net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6944_ _0517_ clknet_leaf_60_core_clock dmmu1.page_table\[2\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_46_1602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6875_ _0448_ clknet_leaf_66_core_clock dmmu1.page_table\[7\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5826_ _1976_ _2484_ _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__3287__B _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5573__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5757_ _2775_ _0391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input382_I ic1_wb_stb vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4708_ _2105_ _2138_ _2141_ immu_1.page_table\[10\]\[10\] _2153_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5688_ _2101_ _2726_ _2728_ net905 _2737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input76_I c0_sr_bus_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4128__A2 net230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4639_ _2113_ _0744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3887__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3431__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6309_ _0691_ clknet_leaf_96_core_clock immu_1.page_table\[3\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5089__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5628__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3639__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6053__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4064__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5261__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5800__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3811__A1 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_3_3_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6697__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5013__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3197__B _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4367__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_5_core_clock_I clknet_4_1__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7183__I net402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_2044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3422__S0 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_2303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4827__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput260 dcache_wb_o_dat[13] net260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput271 dcache_wb_o_dat[9] net271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput282 ic0_mem_data[14] net282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput293 ic0_mem_data[24] net293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4055__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4990_ net103 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_58_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3102__I0 net133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3941_ _1408_ _1599_ _1604_ _1605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_19_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3872_ immu_1.page_table\[0\]\[5\] immu_1.page_table\[1\]\[5\] immu_1.page_table\[2\]\[5\]
+ immu_1.page_table\[3\]\[5\] _1435_ _1469_ _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6660_ _0233_ clknet_leaf_15_core_clock dmmu0.page_table\[11\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5611_ _2693_ _0327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5555__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5555__B2 dmmu0.page_table\[3\]\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6591_ _0164_ clknet_leaf_8_core_clock immu_0.page_table\[3\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5542_ _2654_ _0297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5307__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ _2444_ _2613_ _2615_ dmmu0.page_table\[4\]\[0\] _2616_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput701 net701 inner_wb_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3318__B1 _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4424_ _1981_ _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_22_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4355_ _1866_ _1927_ _1929_ net1055 _1938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7143_ net398 net613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3126__I _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3306_ net158 _0893_ _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7074_ net358 net511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4286_ _1890_ _1894_ _1897_ _1898_ _0606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4818__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_2051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3237_ _0982_ _0983_ _0842_ _0984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6025_ _2792_ _2924_ _2926_ dmmu1.page_table\[3\]\[6\] _2933_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input130_I c1_o_mem_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5491__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_2095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input228_I dcache_mem_o_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3168_ dmmu1.page_table\[8\]\[0\] dmmu1.page_table\[9\]\[0\] dmmu1.page_table\[10\]\[0\]
+ dmmu1.page_table\[11\]\[0\] _0899_ _0902_ _0918_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_55_1203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6035__A2 _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3099_ _0852_ net539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4046__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_82_core_clock_I clknet_4_10__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4597__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5794__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6927_ _0500_ clknet_leaf_59_core_clock dmmu1.page_table\[3\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3729__C _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6858_ _0431_ clknet_leaf_50_core_clock dmmu1.page_table\[8\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5809_ _2809_ _0409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_1832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4349__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6789_ _0362_ clknet_leaf_43_core_clock dmmu1.page_table\[13\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3404__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output447_I net447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4521__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3955__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4037__A1 net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5234__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7178__I net397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_2010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3260__A2 dmmu1.page_table\[14\]\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3563__A3 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6712__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4140_ net86 _1786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4071_ _1726_ _1729_ _1731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6862__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5473__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6017__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4579__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4973_ _2318_ _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_58_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6712_ _0285_ clknet_leaf_29_core_clock dmmu0.page_table\[13\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3924_ immu_0.page_table\[12\]\[6\] immu_0.page_table\[13\]\[6\] immu_0.page_table\[14\]\[6\]
+ immu_0.page_table\[15\]\[6\] _1424_ _1455_ _1588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_74_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6643_ _0216_ clknet_leaf_30_core_clock dmmu0.page_table\[15\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3855_ _1517_ _1520_ _1440_ _1521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_0_27_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6242__CLK clknet_leaf_85_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3786_ _1454_ net664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6574_ _0147_ clknet_leaf_21_core_clock immu_0.page_table\[4\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5525_ net94 _2629_ _2631_ net752 _2644_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4751__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input178_I c1_o_req_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3284__C _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput520 net520 dcache_mem_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5456_ _2605_ _0260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6392__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput531 net531 dcache_mem_addr[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_30_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput542 net542 dcache_mem_cache_enable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput553 net553 dcache_mem_i_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4407_ _1866_ _1957_ _1959_ net873 _1968_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput564 net564 dcache_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5700__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput575 net575 dcache_wb_i_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5387_ _2564_ _0232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput586 net586 ic0_mem_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_61_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input345_I ic1_mem_data[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7126_ net71 net594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput597 net597 ic0_mem_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4338_ _1928_ _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_10_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input39_I c0_o_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7057_ net294 net445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4269_ _1864_ _1876_ _1878_ net899 _1886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4267__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6008_ _2922_ _0495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4019__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3242__A2 _0979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3873__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5519__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3475__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output564_I net564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6885__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6265__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_13__f_core_clock clknet_3_6_0_core_clock clknet_4_13__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_83_2697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3864__S0 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3784__A3 _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3640_ _1323_ net690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3571_ net222 _1204_ _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_24_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5310_ _2520_ _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6290_ _0672_ clknet_leaf_101_core_clock dmmu0.page_table\[0\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5241_ _2479_ _0171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3919__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4497__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4041__S0 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3544__I0 net149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5172_ _2269_ _2430_ _2432_ net1064 _2436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4123_ _1773_ net466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput2 c0_o_c_instr_long net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4054_ immu_0.page_table\[4\]\[10\] immu_0.page_table\[5\]\[10\] immu_0.page_table\[6\]\[10\]
+ immu_0.page_table\[7\]\[10\] _1370_ _1391_ _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5997__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6608__CLK clknet_leaf_24_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4235__I net207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3279__C _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _2275_ _2299_ _2302_ net1083 _2309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_1072 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6758__CLK clknet_leaf_99_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3907_ _1570_ _1571_ _1366_ _1572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4972__A2 _2316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4887_ _2260_ _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_62_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input295_I ic0_mem_data[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6626_ _0199_ clknet_leaf_29_core_clock dmmu0.page_table\[12\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3838_ _1440_ _1504_ _1505_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6557_ _0130_ clknet_leaf_21_core_clock immu_0.page_table\[6\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5921__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3769_ _1437_ _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_30_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5508_ _2635_ _0282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6488_ _0061_ clknet_leaf_13_core_clock dmmu0.page_table\[7\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5439_ _2594_ _0254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3515__S _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7109_ net400 net577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6288__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4660__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output681_I net681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6165__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_19_core_clock_I clknet_4_4__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7191__I net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A1 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_29_Left_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5676__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_72_2387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5428__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__A1 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_85_2759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_30_core_clock clknet_4_5__leaf_core_clock clknet_leaf_30_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_76_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6900__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Left_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4810_ _1809_ _2208_ _2210_ immu_0.page_table\[13\]\[5\] _2216_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_1971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4403__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5790_ _2105_ _2777_ _2779_ dmmu1.page_table\[10\]\[10\] _2798_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5600__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3837__S0 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4741_ _1790_ _2173_ _2174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_22_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4954__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4672_ _2067_ _2123_ _2125_ net1032 _2132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_12_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6411_ _0793_ clknet_leaf_112_core_clock immu_0.page_table\[14\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_42_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5903__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3623_ _1308_ net268 _1315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4706__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6342_ _0724_ clknet_leaf_77_core_clock immu_1.page_table\[14\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3554_ net139 net34 _1267_ _1277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_47_Left_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6273_ _0655_ clknet_leaf_90_core_clock immu_1.page_table\[6\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3485_ dmmu0.page_table\[4\]\[11\] dmmu0.page_table\[5\]\[11\] dmmu0.page_table\[6\]\[11\]
+ dmmu0.page_table\[7\]\[11\] _0864_ _0867_ _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_62_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5224_ _1789_ _2468_ _2469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_55_1862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_51_1737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3134__I _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5155_ _2328_ _2414_ _2416_ net1095 _2425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4890__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3693__A2 net311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4106_ _1350_ net327 _1360_ _1762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5086_ _2385_ _0110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_32_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4037_ net9 immu_0.high_addr_off\[4\] _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_21_core_clock_I clknet_4_4__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input210_I c1_sr_bus_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4642__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_56_Left_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input308_I ic0_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5988_ _2912_ _0485_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4939_ _1977_ _2297_ _2298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_19_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6147__A1 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6609_ _0182_ clknet_leaf_15_core_clock immu_0.page_table\[1\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_65_Left_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5370__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3220__I2 dmmu1.page_table\[14\]\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3381__A1 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3133__A1 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output527_I net527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3044__I _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3684__A2 net324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6923__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6083__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_74_Left_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5830__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5189__A2 _1971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3819__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_2055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4397__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7186__I net390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4149__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_2552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5897__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_74_2427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_2438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_2075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_2449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3372__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6453__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3382__C _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3270_ _1014_ _0858_ _1015_ _1016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4321__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4872__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6960_ _0533_ clknet_leaf_65_core_clock dmmu1.page_table\[1\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_1058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5911_ _2849_ _2856_ _2858_ net836 _2868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_2019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6891_ _0464_ clknet_leaf_61_core_clock dmmu1.page_table\[6\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_1318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5842_ _1811_ _2819_ _2821_ dmmu0.page_table\[1\]\[6\] _2828_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_87_core_clock_I clknet_4_10__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5773_ _2787_ _0395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4927__A2 _2285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_20_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4724_ _1806_ _2157_ _2159_ net896 _2164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6129__A1 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4655_ _2121_ _0752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3129__I _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3606_ _0814_ net328 net659 _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput60 c0_o_req_addr[10] net60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput71 c0_o_req_addr[6] net71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5352__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput82 c0_sr_bus_addr[15] net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4586_ _2081_ _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_57_1924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput93 c0_sr_bus_data_o[10] net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_57_1935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6325_ _0707_ clknet_leaf_70_core_clock dmmu1.page_table\[14\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3537_ _1268_ net554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_1594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input160_I c1_o_mem_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input258_I dcache_wb_o_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6256_ _0638_ clknet_leaf_95_core_clock immu_1.page_table\[5\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3468_ dmmu1.page_table\[8\]\[11\] dmmu1.page_table\[9\]\[11\] dmmu1.page_table\[10\]\[11\]
+ dmmu1.page_table\[11\]\[11\] _0898_ _0901_ _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__6946__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5207_ _2458_ _0158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6187_ net738 _3025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3399_ net48 dmmu0.long_off_reg\[3\] _1140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_4_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3666__A2 net320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5138_ _2415_ _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_77_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input21_I c0_o_mem_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ _2273_ _2367_ _2369_ immu_0.page_table\[8\]\[5\] _2375_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4615__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5812__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6326__CLK clknet_leaf_70_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4379__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5455__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6476__CLK clknet_leaf_92_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3106__A1 net50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4303__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3657__A2 net318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3930__C _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_2220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_2242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_63_2106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_63_2117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_2017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5031__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6819__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3593__A1 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4790__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4440_ _1990_ _0668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5334__A2 _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold107 immu_0.page_table\[3\]\[1\] net841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold118 dmmu0.page_table\[9\]\[9\] net852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold129 immu_1.page_table\[11\]\[8\] net863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3345__A1 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4371_ _1852_ _1942_ _1944_ net1050 _1948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6110_ _2981_ _0538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_1024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3322_ dmmu1.page_table\[12\]\[6\] dmmu1.page_table\[13\]\[6\] dmmu1.page_table\[14\]\[6\]
+ dmmu1.page_table\[15\]\[6\] _0888_ _0901_ _1066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7090_ net344 net497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4001__C _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6041_ _1770_ _2940_ _2942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_33_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3253_ _0931_ _0995_ _0998_ _0896_ _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_20_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3648__A2 net370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4845__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3184_ net106 _0932_ _0933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__6047__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4508__I _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6349__CLK clknet_leaf_62_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6943_ _0516_ clknet_leaf_60_core_clock dmmu1.page_table\[2\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_46_1603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6874_ _0447_ clknet_leaf_55_core_clock dmmu1.page_table\[7\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5825_ _2817_ _0417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6499__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5756_ _2049_ _2759_ _2761_ net884 _2775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5573__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4707_ _2152_ _0773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5687_ _2736_ _0360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input375_I ic1_wb_adr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4638_ _2059_ _2108_ _2110_ immu_1.page_table\[12\]\[2\] _2113_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input69_I c0_o_req_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4569_ _1866_ _2053_ _2055_ net849 _2071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3887__A2 _1546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3431__S1 _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6308_ _0690_ clknet_leaf_89_core_clock immu_1.page_table\[3\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5089__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6239_ _0621_ clknet_leaf_82_core_clock immu_1.page_table\[2\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3639__A2 net261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3523__S _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3195__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4064__A2 _1723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5261__A1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output594_I net594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5013__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3575__A1 net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4772__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_2012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3327__A1 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4102__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3422__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4827__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3433__S _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput250 dcache_wb_adr[5] net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput261 dcache_wb_o_dat[14] net261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6029__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput272 dcache_wb_sel[0] net272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput283 ic0_mem_data[15] net283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput294 ic0_mem_data[25] net294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_1006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3102__I1 net28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6641__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3940_ _1446_ _1601_ _1603_ _1604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_74_905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3871_ _1306_ _1523_ _1534_ _1536_ net667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_6_1282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5610_ _2527_ _2681_ _2684_ net803 _2693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5555__A2 _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6590_ _0163_ clknet_leaf_19_core_clock immu_0.page_table\[3\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6791__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4763__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5541_ _2457_ _2647_ _2649_ dmmu0.page_table\[3\]\[4\] _2654_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5307__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5472_ _2614_ _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_67_1878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3318__A1 _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput702 net702 inner_wb_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4515__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4423_ _1980_ _1978_ _1981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3318__B2 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7142_ net397 net612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4354_ _1937_ _0635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_6_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3305_ net150 dmmu1.long_off_reg\[0\] _1050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7073_ net357 net510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4285_ net736 _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3343__S _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4818__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6024_ _2932_ _0501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3236_ _0915_ _0895_ _0983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5491__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3167_ _0897_ _0916_ _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input123_I c1_o_mem_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3098_ net131 net26 _0850_ _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4046__A2 net244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6926_ _0499_ clknet_leaf_54_core_clock dmmu1.page_table\[3\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ _0430_ clknet_leaf_101_core_clock dmmu0.page_table\[1\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5808_ _2788_ _2802_ _2804_ dmmu1.page_table\[9\]\[4\] _2809_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6788_ _0361_ clknet_leaf_45_core_clock dmmu1.page_table\[13\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5739_ _2766_ _0382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3309__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3404__S1 _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6514__CLK clknet_leaf_2_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3168__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_1440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6664__CLK clknet_leaf_109_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3052__I _0826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5234__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3096__I0 net130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3796__A1 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5537__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6194__CLK clknet_leaf_2_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5170__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4070_ _1726_ _1729_ _1730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5473__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_2034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3087__I0 net126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4972_ _2300_ _2316_ _2318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_clkbuf_leaf_26_core_clock_I clknet_4_5__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6711_ _0284_ clknet_leaf_33_core_clock dmmu0.page_table\[13\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_1388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3331__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4984__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3923_ _1383_ _1584_ _1586_ _1587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_15_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6642_ _0215_ clknet_leaf_32_core_clock dmmu0.page_table\[15\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3854_ _1518_ _1519_ _1446_ _1520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6573_ _0146_ clknet_leaf_27_core_clock immu_0.page_table\[4\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3785_ net235 _1453_ _1360_ _1454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5524_ _2643_ _0290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6537__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5455_ immu_1.high_addr_off\[1\] _1846_ _2603_ _2605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_2051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput510 net510 c1_i_req_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3137__I _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput521 net521 dcache_mem_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput532 net532 dcache_mem_addr[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput543 net543 dcache_mem_i_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4406_ _1967_ _0657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput554 net554 dcache_mem_i_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5386_ _2527_ _2553_ _2555_ dmmu0.page_table\[11\]\[8\] _2564_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput565 net565 dcache_wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput576 net576 dcache_wb_i_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3711__A1 net385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7125_ net70 net593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput587 net587 ic0_mem_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput598 net598 ic0_mem_cache_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4337_ _1912_ _1926_ _1928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6687__CLK clknet_leaf_91_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input240_I dcache_wb_adr[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input338_I ic1_mem_data[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7056_ net293 net444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4268_ _1885_ _0601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4267__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6007_ net200 _2906_ _2908_ dmmu1.page_table\[4\]\[12\] _2922_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3219_ dmmu1.page_table\[4\]\[2\] dmmu1.page_table\[5\]\[2\] dmmu1.page_table\[6\]\[2\]
+ dmmu1.page_table\[7\]\[2\] _0889_ _0931_ _0967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_4199_ _1830_ net196 _1833_ _1834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_59_1170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_2__f_core_clock clknet_3_1_0_core_clock clknet_4_2__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4019__A2 net243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_2011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3600__I _1300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_1490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3778__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3322__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6909_ _0482_ clknet_leaf_64_core_clock dmmu1.page_table\[5\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_1928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3873__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5519__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5463__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold290 immu_1.page_table\[5\]\[7\] net1024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_79_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_20_core_clock clknet_4_4__leaf_core_clock clknet_leaf_20_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_1877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7189__I net393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_2698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3864__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3666__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4718__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_1940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4194__A1 _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3570_ _1285_ net418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3941__A1 _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5143__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5240_ _2461_ _2470_ _2472_ immu_0.page_table\[2\]\[6\] _2479_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4497__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4041__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5694__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3544__I1 net44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Right_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5171_ _2435_ _0145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4122_ net212 _0831_ _1773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5446__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4249__A2 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4053_ _1708_ _1711_ _1579_ _1713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_56_2033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput3 c0_o_c_instr_page net3 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5997__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_2017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4955_ _2308_ _0056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_27_Right_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3906_ _1396_ immu_0.page_table\[9\]\[5\] _1390_ _1571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4886_ _1977_ _2259_ _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6625_ _0198_ clknet_leaf_29_core_clock dmmu0.page_table\[12\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3837_ immu_1.page_table\[8\]\[3\] immu_1.page_table\[9\]\[3\] immu_1.page_table\[10\]\[3\]
+ immu_1.page_table\[11\]\[3\] _1474_ _1469_ _1504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_15_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input190_I c1_sr_bus_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input288_I ic0_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5382__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6556_ _0129_ clknet_leaf_23_core_clock immu_0.page_table\[6\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3768_ _1434_ _1436_ net705 _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5507_ _2453_ _2630_ _2632_ dmmu0.page_table\[13\]\[2\] _2635_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3932__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6487_ _0060_ clknet_leaf_13_core_clock dmmu0.page_table\[7\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3699_ net312 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_63_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5438_ _2529_ _2582_ _2584_ net881 _2594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_36_Right_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input51_I c0_o_mem_high_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5082__I _2381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5369_ _2554_ _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7108_ net399 net576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_94_core_clock_I clknet_4_8__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7039_ net306 net457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3531__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3999__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4660__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6702__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4948__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_2104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6852__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3923__A1 _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Right_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_76_2491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_2000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4479__A2 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5676__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_2388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5428__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6232__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5979__A2 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Right_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6382__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5600__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4403__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3837__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4740_ _2154_ _2172_ _2173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_51_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4671_ _2131_ _0758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6410_ _0792_ clknet_leaf_0_core_clock immu_0.page_table\[14\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3622_ _1314_ net696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_42_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5903__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_72_Right_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_12_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3914__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ _0723_ clknet_leaf_73_core_clock immu_1.page_table\[14\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3553_ _1276_ net547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5116__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6272_ _0654_ clknet_leaf_85_core_clock immu_1.page_table\[6\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3843__C _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3484_ _0877_ _1220_ _1222_ _0958_ _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_42_1910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5223_ _1971_ _2172_ _2468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5154_ _2424_ _0139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_36_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4890__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4105_ _1348_ net381 _1761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5085_ _2258_ _2382_ _2384_ net847 _2385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_81_Right_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4036_ net9 immu_0.high_addr_off\[4\] _1697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6725__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4642__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3150__I net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input203_I c1_sr_bus_data_o[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_1678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5987_ _2784_ _2907_ _2909_ net988 _2912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6875__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4938_ _1780_ _2296_ _2297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_19_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input99_I c0_sr_bus_data_o[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_30 net397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6147__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4869_ _2250_ _0028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6608_ _0181_ clknet_leaf_24_core_clock immu_0.page_table\[1\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3905__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6539_ _0112_ clknet_leaf_6_core_clock immu_0.page_table\[7\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_7__f_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6255__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6083__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3516__S0 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_2094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4156__I _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5830__A1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_2170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_2034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3819__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4397__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_2045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_2056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5594__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4149__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5346__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5897__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_2428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_2439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4321__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4872__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6898__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5910_ _2867_ _0452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6890_ _0463_ clknet_leaf_56_core_clock dmmu1.page_table\[6\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5841_ _2827_ _0423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5772_ _2786_ _2778_ _2780_ net1089 _2787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_44_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__B1 _2665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4723_ _2163_ _0778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_40_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6129__A2 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4654_ _2105_ _2107_ _2109_ net1001 _2121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput50 c0_o_mem_high_addr[5] net50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3605_ _1304_ net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6278__CLK clknet_leaf_95_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput61 c0_o_req_addr[11] net61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput72 c0_o_req_addr[7] net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4585_ _2061_ _2075_ _2077_ immu_1.page_table\[14\]\[3\] _2081_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_57_1914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput83 c0_sr_bus_addr[1] net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_57_1925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput94 c0_sr_bus_data_o[11] net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6324_ _0706_ clknet_leaf_70_core_clock dmmu1.page_table\[14\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_1936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3994__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3536_ net145 net40 _1267_ _1268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6255_ _0637_ clknet_leaf_86_core_clock immu_1.page_table\[5\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3467_ _0897_ _1205_ _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input153_I c1_o_mem_high_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5206_ _2457_ _2447_ _2449_ immu_0.page_table\[3\]\[4\] _2458_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6186_ _3024_ _0571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3398_ _1118_ _1124_ _1139_ net528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_4_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5137_ _1980_ _2413_ _2415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3081__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input320_I ic0_wb_adr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6065__A1 net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5068_ _2374_ _0103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5812__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input14_I c0_o_mem_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4615__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4019_ net659 net243 _1681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4091__A3 _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Right_0 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4379__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3051__A1 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_1176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3106__A2 net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4303__A1 net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4854__A2 _2240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_2221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5654__I1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4082__A3 _1741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3290__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5406__I1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_14_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6420__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5319__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4790__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3593__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold108 immu_0.page_table\[14\]\[0\] net842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold119 dmmu0.page_table\[12\]\[1\] net853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4542__A1 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4370_ _1947_ _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6570__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3321_ dmmu1.page_table\[0\]\[6\] dmmu1.page_table\[1\]\[6\] dmmu1.page_table\[2\]\[6\]
+ dmmu1.page_table\[3\]\[6\] _0888_ _0910_ _1065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_10_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6040_ _2940_ _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3252_ _0889_ _0996_ _0997_ _0902_ _0998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_28_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I c0_o_instr_long_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4845__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3183_ net158 _0932_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_59_1522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6047__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6942_ _0515_ clknet_leaf_58_core_clock dmmu1.page_table\[2\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_1604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6873_ _0446_ clknet_leaf_52_core_clock dmmu1.page_table\[7\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5824_ _2049_ _2801_ _2803_ net1060 _2817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5755_ _2774_ _0390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4706_ _2103_ _2139_ _2142_ net829 _2152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5686_ _2069_ _2726_ _2728_ dmmu1.page_table\[13\]\[7\] _2736_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6913__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4637_ _2112_ _0743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_66_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input270_I dcache_wb_o_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4533__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3336__A2 _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input368_I ic1_wb_adr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4568_ _2070_ _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_33_core_clock_I clknet_4_7__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6307_ _0689_ clknet_leaf_83_core_clock immu_1.page_table\[3\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3519_ _0896_ _1256_ _1257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _1866_ _2014_ _2016_ immu_1.page_table\[3\]\[8\] _2025_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3804__S _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5089__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6238_ _0620_ clknet_leaf_91_core_clock immu_1.page_table\[2\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4297__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6169_ _2029_ _2601_ _3015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3195__S1 _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3895__I0 _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5261__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6443__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5549__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5013__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_1659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_2051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output587_I net587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4221__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3575__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6593__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3327__A2 _1068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3958__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4827__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput240 dcache_wb_adr[18] net240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput251 dcache_wb_adr[6] net251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6029__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput262 dcache_wb_o_dat[15] net262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput273 dcache_wb_sel[1] net273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput284 ic0_mem_data[16] net284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput295 ic0_mem_data[26] net295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5788__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3263__A1 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3870_ _1535_ net238 _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6936__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4763__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5540_ _2653_ _0296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_82_972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5471_ _2300_ _2612_ _2614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_48_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput703 net703 inner_wb_stb vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4515__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4422_ _1769_ _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_2_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4515__B2 dmmu1.page_table\[14\]\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5712__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7141_ net396 net611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4353_ _1864_ _1927_ _1929_ net1024 _1937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_6_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3304_ _0915_ _1042_ _1044_ _1046_ _1048_ _1049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_7072_ net356 net509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4284_ _1896_ _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6316__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4818__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6023_ _2790_ _2924_ _2926_ dmmu1.page_table\[3\]\[5\] _2932_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3235_ _0980_ _0981_ _0907_ _0982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_99_core_clock_I clknet_4_3__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5491__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_2097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3166_ dmmu1.page_table\[12\]\[0\] dmmu1.page_table\[13\]\[0\] dmmu1.page_table\[14\]\[0\]
+ dmmu1.page_table\[15\]\[0\] _0899_ _0902_ _0916_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_55_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6466__CLK clknet_leaf_32_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3097_ _0851_ net538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input116_I c1_o_instr_long_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6925_ _0498_ clknet_leaf_53_core_clock dmmu1.page_table\[3\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6856_ _0429_ clknet_leaf_100_core_clock dmmu0.page_table\[1\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5807_ _2808_ _0408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_1968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3999_ _1434_ _1660_ _1661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6787_ _0360_ clknet_leaf_44_core_clock dmmu1.page_table\[13\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5738_ _2061_ _2760_ _2762_ net1088 _2766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input81_I c0_sr_bus_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5669_ _2725_ _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_27_1318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3168__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6809__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_2017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_10_core_clock clknet_4_3__leaf_core_clock clknet_leaf_10_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3493__A1 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4690__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output502_I net502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5234__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6959__CLK clknet_leaf_64_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3096__I1 net25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4164__I _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4745__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6339__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5170__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6489__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5473__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3484__A1 _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_99_core_clock clknet_4_3__leaf_core_clock clknet_leaf_99_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3236__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4971_ _2316_ _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3087__I1 net21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4433__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6710_ _0283_ clknet_leaf_29_core_clock dmmu0.page_table\[13\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4984__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3922_ _1368_ _1585_ _1586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3331__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4984__B2 dmmu0.page_table\[14\]\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6641_ _0214_ clknet_leaf_29_core_clock dmmu0.page_table\[15\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3853_ immu_1.page_table\[0\]\[4\] immu_1.page_table\[1\]\[4\] immu_1.page_table\[2\]\[4\]
+ immu_1.page_table\[3\]\[4\] _1409_ _1442_ _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_41_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4736__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5933__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3784_ _1422_ _1427_ _1432_ _1452_ _1453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_6572_ _0145_ clknet_leaf_20_core_clock immu_0.page_table\[4\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5523_ _2531_ _2629_ _2631_ net991 _2643_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5454_ _2604_ _0259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput500 net500 c1_i_req_data[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput511 net511 c1_i_req_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput522 net522 dcache_mem_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4405_ _1864_ _1957_ _1959_ net769 _1967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput533 net533 dcache_mem_addr[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5161__A1 _1972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput544 net544 dcache_mem_i_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5385_ _2563_ _0231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput555 net555 dcache_mem_i_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput566 net566 dcache_wb_i_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput577 net577 dcache_wb_i_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3172__B1 _0921_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7124_ net69 net592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4336_ _1926_ _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput588 net588 ic0_mem_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput599 net599 ic0_mem_ppl_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_5_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7055_ net292 net443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4267_ _1861_ _1876_ _1878_ immu_1.page_table\[7\]\[6\] _1885_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input233_I dcache_wb_adr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6006_ _2921_ _0494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3218_ _0964_ _0965_ _0842_ _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_1761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4198_ _1831_ _1832_ _1833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4672__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3149_ _0898_ _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_2050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input400_I inner_wb_i_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3227__A1 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6908_ _0481_ clknet_leaf_65_core_clock dmmu1.page_table\[5\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3322__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6839_ _0412_ clknet_leaf_45_core_clock dmmu1.page_table\[9\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3529__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output452_I net452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6631__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold280 dmmu1.page_table\[8\]\[1\] net1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold291 dmmu0.page_table\[12\]\[6\] net1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4159__I net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6781__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4966__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_2699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4718__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4194__A2 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5654__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5143__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5694__A2 _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5170_ _2267_ _2430_ _2432_ net1038 _2435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4121_ _1306_ _1302_ _0816_ net641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_78_1024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__A2 net379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4052_ _1708_ _1711_ _1712_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3457__A1 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 c0_o_icache_flush net4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_1934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4954_ _2273_ _2299_ _2302_ dmmu0.page_table\[7\]\[5\] _2308_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3905_ _1385_ immu_0.page_table\[8\]\[5\] _1570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6159__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ _1779_ _1972_ _2259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_15_1096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6624_ _0197_ clknet_leaf_12_core_clock immu_0.page_table\[0\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3836_ _1408_ _1501_ _1502_ _1503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_46_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5382__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3767_ immu_1.page_table\[0\]\[1\] immu_1.page_table\[1\]\[1\] immu_1.page_table\[8\]\[1\]
+ immu_1.page_table\[9\]\[1\] _1435_ _1415_ _1436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6555_ _0128_ clknet_leaf_22_core_clock immu_0.page_table\[6\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3148__I _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6654__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input183_I c1_sr_bus_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5506_ _2634_ _0281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6486_ _0059_ clknet_leaf_36_core_clock dmmu0.page_table\[7\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3698_ _1367_ _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_63_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5437_ _2593_ _0253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input350_I ic1_mem_data[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5368_ _2300_ _2552_ _2554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4893__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input44_I c0_o_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7107_ net398 net575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4319_ _1852_ _1911_ _1914_ net919 _1918_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5299_ net104 _2502_ _2504_ immu_0.page_table\[0\]\[9\] _2513_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7038_ net305 net456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3448__A1 net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_2_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4948__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_76_2492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_0_core_clock clknet_4_0__leaf_core_clock clknet_leaf_0_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4479__A3 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5676__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3687__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_107_core_clock clknet_4_2__leaf_core_clock clknet_leaf_107_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_24_1877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5428__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3439__A1 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4636__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__A3 _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_2049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_2073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5061__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3298__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5600__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3611__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6677__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4670_ _2065_ _2123_ _2125_ net1084 _2131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3621_ _1308_ net267 _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_42_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5364__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3552_ net138 net33 _1267_ _1276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6340_ _0722_ clknet_leaf_73_core_clock immu_1.page_table\[14\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6271_ _0653_ clknet_leaf_91_core_clock immu_1.page_table\[6\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5116__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3483_ _0875_ _1221_ _1222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5222_ _2467_ _0164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_1343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_core_clock_I clknet_4_6__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5153_ _2277_ _2414_ _2416_ net1022 _2424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_36_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4104_ _1758_ _1759_ _1760_ net701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5084_ _2383_ _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_58_1417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4035_ net107 _1685_ _1695_ _1696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_49_1679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5986_ _2911_ _0484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4937_ _1778_ net84 _2296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_34_1483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input398_I inner_wb_i_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_20 net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_31 net397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4868_ _1809_ _2242_ _2244_ net819 _2250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_10_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6607_ _0180_ clknet_leaf_19_core_clock immu_0.page_table\[1\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3819_ immu_0.page_table\[0\]\[3\] immu_0.page_table\[1\]\[3\] immu_0.page_table\[2\]\[3\]
+ immu_0.page_table\[3\]\[3\] _1424_ _1455_ _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_43_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4799_ _2209_ _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_16_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6538_ _0111_ clknet_leaf_3_core_clock immu_0.page_table\[7\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6469_ _0042_ clknet_leaf_16_core_clock dmmu0.page_table\[8\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3669__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3542__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_2051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6083__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3516__S1 net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5291__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5830__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3841__A1 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_2171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5043__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_2182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_40_core_clock_I clknet_4_6__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_2046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5594__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4397__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_2057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4172__I _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5346__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4149__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5897__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_2429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4321__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4609__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4085__A1 net11 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5282__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ _1808_ _2819_ _2821_ net1091 _2827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5585__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5771_ _1851_ _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_12_1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3200__B _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4722_ _1803_ _2157_ _2159_ immu_0.page_table\[15\]\[3\] _2163_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4653_ _2120_ _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput40 c0_o_mem_data[5] net40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3604_ inner_wb_arbiter.o_sel_sig _1304_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
Xinput51 c0_o_mem_high_addr[6] net51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput62 c0_o_req_addr[12] net62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3899__A1 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4584_ _2080_ _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput73 c0_o_req_addr[8] net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_57_1915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput84 c0_sr_bus_addr[2] net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput95 c0_sr_bus_data_o[12] net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6323_ _0705_ clknet_leaf_70_core_clock dmmu1.page_table\[14\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_1926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3535_ _0840_ _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_29_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3994__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6254_ _0636_ clknet_leaf_87_core_clock immu_1.page_table\[5\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3466_ dmmu1.page_table\[12\]\[11\] dmmu1.page_table\[13\]\[11\] dmmu1.page_table\[14\]\[11\]
+ dmmu1.page_table\[15\]\[11\] _0898_ _0901_ _1205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_38_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ _1805_ _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6185_ dmmu1.long_off_reg\[7\] _1864_ _3016_ _3024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3397_ net106 net158 _0884_ _1138_ _1139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_42_1796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input146_I c1_o_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5136_ _2413_ _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_4_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6065__A2 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5067_ _2271_ _2367_ _2369_ net747 _2374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5273__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6842__CLK clknet_leaf_67_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input313_I ic0_wb_adr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5812__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4018_ _1654_ _1664_ _1669_ _1679_ _1680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_7_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3823__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5025__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4379__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6992__CLK clknet_leaf_94_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5969_ _2847_ _2890_ _2892_ net1096 _2901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3051__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4000__A1 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3434__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4839__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output532_I net532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3106__A3 net52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4303__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput400 inner_wb_i_dat[5] net400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_76_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_2222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4067__A1 net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_2233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3814__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_2119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5567__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3042__A2 net559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5319__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4790__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6715__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold109 dmmu1.page_table\[12\]\[2\] net843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4542__A2 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5662__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3320_ dmmu1.page_table\[4\]\[6\] dmmu1.page_table\[5\]\[6\] dmmu1.page_table\[6\]\[6\]
+ dmmu1.page_table\[7\]\[6\] _0888_ _0910_ _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_21_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3750__B1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3251_ _0908_ dmmu1.page_table\[0\]\[4\] _0997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_33_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6865__CLK clknet_leaf_46_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3182_ _0901_ _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_20_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6047__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4058__A1 _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5255__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6941_ _0514_ clknet_leaf_58_core_clock dmmu1.page_table\[2\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3805__A1 _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_1605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6872_ _0445_ clknet_leaf_55_core_clock dmmu1.page_table\[7\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5007__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5823_ _2816_ _0416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6245__CLK clknet_leaf_94_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_1420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5754_ _2047_ _2759_ _2761_ net894 _2774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3865__B _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4705_ _2151_ _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5685_ _2735_ _0359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4636_ _2057_ _2108_ _2110_ net750 _2112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5730__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4567_ _2069_ _2053_ _2055_ net765 _2070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3156__I _0905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input263_I dcache_wb_o_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6306_ _0688_ clknet_leaf_91_core_clock immu_1.page_table\[3\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3518_ dmmu1.page_table\[12\]\[12\] dmmu1.page_table\[13\]\[12\] dmmu1.page_table\[14\]\[12\]
+ dmmu1.page_table\[15\]\[12\] _0886_ net121 _1256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4498_ _2024_ _0692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_1137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6237_ _0619_ clknet_leaf_95_core_clock immu_1.page_table\[2\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3449_ net154 dmmu1.long_off_reg\[4\] _1189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4297__A1 _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6168_ _1764_ _1767_ _3014_ _0563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5119_ _2404_ _0124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4049__A1 net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6099_ _1891_ _1892_ _2030_ _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__5246__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5549__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4221__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6738__CLK clknet_leaf_46_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4772__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4450__I net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3407__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3958__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6888__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5485__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput230 dcache_wb_4_burst net230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput241 dcache_wb_adr[19] net241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput252 dcache_wb_adr[7] net252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6029__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput263 dcache_wb_o_dat[1] net263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput274 dcache_wb_stb net274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput285 ic0_mem_data[17] net285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput296 ic0_mem_data[27] net296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_89_core_clock clknet_4_8__leaf_core_clock clknet_leaf_89_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5788__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3894__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4763__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5470_ _2612_ _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_48_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4421_ _1978_ _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput704 net704 inner_wb_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4515__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5712__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7140_ net389 net604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4352_ _1936_ _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_1435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3303_ _0897_ _1047_ _0912_ _1048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_22_1419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7071_ net353 net506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4283_ _1895_ _1893_ _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5191__I _2446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3234_ dmmu1.page_table\[0\]\[3\] dmmu1.page_table\[1\]\[3\] dmmu1.page_table\[2\]\[3\]
+ dmmu1.page_table\[3\]\[3\] _0899_ _0902_ _0981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_59_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6022_ _2931_ _0500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3165_ net123 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5228__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3096_ net130 net25 _0850_ _0851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4535__I net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6924_ _0497_ clknet_leaf_56_core_clock dmmu1.page_table\[3\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4451__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input109_I c1_o_icache_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6855_ _0428_ clknet_leaf_100_core_clock dmmu0.page_table\[1\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5806_ _2786_ _2802_ _2804_ net935 _2808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_1971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4203__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6786_ _0359_ clknet_leaf_46_core_clock dmmu1.page_table\[13\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3998_ immu_1.page_table\[12\]\[8\] immu_1.page_table\[13\]\[8\] immu_1.page_table\[14\]\[8\]
+ immu_1.page_table\[15\]\[8\] _1441_ _1540_ _1660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_73_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5737_ _2765_ _0381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5951__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3087__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input380_I ic1_wb_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_2009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5668_ _1828_ _2028_ _2031_ _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_5_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input74_I c0_o_req_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4619_ _2069_ _2090_ _2092_ net844 _2100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_1379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5599_ _2687_ _0321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6410__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3550__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5219__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3493__A2 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4690__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3876__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6560__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3556__I0 net140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5170__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3181__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6903__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _1977_ _2173_ _2316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__3236__A2 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4433__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5630__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3921_ immu_0.page_table\[0\]\[6\] immu_0.page_table\[1\]\[6\] immu_0.page_table\[2\]\[6\]
+ immu_0.page_table\[3\]\[6\] _1424_ _1455_ _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_50_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4984__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6640_ _0213_ clknet_leaf_30_core_clock dmmu0.page_table\[15\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3852_ immu_1.page_table\[8\]\[4\] immu_1.page_table\[9\]\[4\] immu_1.page_table\[10\]\[4\]
+ immu_1.page_table\[11\]\[4\] _1409_ _1442_ _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__5933__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4736__A2 _2156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6571_ _0144_ clknet_leaf_9_core_clock immu_0.page_table\[4\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3783_ _1433_ _1438_ _1451_ _0813_ _1452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_54_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5522_ _2642_ _0289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5453_ immu_1.high_addr_off\[0\] _1824_ _2603_ _2604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_1688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput501 net501 c1_i_req_data[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4044__S0 _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput512 net512 c1_i_req_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput523 net523 dcache_mem_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_84_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4404_ _1966_ _0656_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput534 net534 dcache_mem_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput545 net545 dcache_mem_i_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5384_ _2463_ _2553_ _2555_ dmmu0.page_table\[11\]\[7\] _2563_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput556 net556 dcache_mem_i_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput567 net567 dcache_wb_i_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3172__B2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7123_ net68 net591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput578 net578 dcache_wb_i_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_5_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4335_ _1828_ _1839_ _1873_ _1926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__3711__A3 net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput589 net589 ic0_mem_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7054_ net291 net442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4266_ _1884_ _0600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6005_ net199 _2906_ _2908_ dmmu1.page_table\[4\]\[11\] _2921_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3217_ _0897_ _0895_ _0965_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3370__S _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4197_ net185 net184 net183 net182 _1832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__4672__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input226_I dcache_mem_o_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6583__CLK clknet_leaf_24_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3148_ _0886_ _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_72_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3079_ _0840_ _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_77_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3227__A2 _0973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3858__S0 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_2057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6907_ _0480_ clknet_leaf_65_core_clock dmmu1.page_table\[5\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6838_ _0411_ clknet_leaf_51_core_clock dmmu1.page_table\[9\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4027__I1 _1687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_45_core_clock_I clknet_4_12__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_1619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6769_ _0342_ clknet_leaf_99_core_clock dmmu0.page_table\[5\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3538__I0 net146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5688__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3163__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold270 dmmu0.page_table\[9\]\[11\] net1004 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_output445_I net445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold281 immu_1.page_table\[6\]\[1\] net1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold292 dmmu1.page_table\[9\]\[8\] net1026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6101__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5860__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4415__A1 _1971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3849__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5612__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4966__A2 _2298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6306__CLK clknet_leaf_91_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4718__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5915__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3963__B _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4026__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6456__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3455__S _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_2__f_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3529__I0 net142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5143__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3154__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4351__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4120_ _1306_ _1302_ _0815_ net640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_23_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4051_ _1699_ _1709_ _1710_ _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__3190__S _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4654__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 c0_o_instr_long_addr[0] net5 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_2035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4953_ _2307_ _0055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3904_ _1391_ _1567_ _1568_ _1569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_30_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3857__C _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6159__A1 _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4884_ _1776_ _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_46_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6623_ _0196_ clknet_leaf_15_core_clock immu_0.page_table\[0\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3835_ _1415_ _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_12_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6554_ _0127_ clknet_leaf_23_core_clock immu_0.page_table\[6\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3766_ _1409_ _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5382__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5505_ _2451_ _2630_ _2632_ net814 _2634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_6_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3393__A1 _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6485_ _0058_ clknet_leaf_32_core_clock dmmu0.page_table\[7\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3697_ _1366_ _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_14_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input176_I c1_o_req_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5436_ _2527_ _2582_ _2584_ dmmu0.page_table\[2\]\[8\] _2593_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6949__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3145__A1 net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5367_ _2552_ _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_1794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input343_I ic1_mem_data[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4893__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7106_ net397 net574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4318_ _1917_ _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5298_ _2512_ _0195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input37_I c0_o_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7037_ net304 net455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4249_ _1872_ net189 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__5842__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_2_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4948__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_1_0_core_clock clknet_0_core_clock clknet_3_1_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_65_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3384__A1 net152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3783__B _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4581__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Left_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4008__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_2493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6173__I1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_2368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_2379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3687__A2 net364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4636__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5061__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3298__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3611__A2 net256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3620_ _1313_ net695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5364__A2 _2535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3693__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3551_ _1275_ net546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6270_ _0652_ clknet_leaf_90_core_clock immu_1.page_table\[6\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5116__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3482_ dmmu0.page_table\[12\]\[11\] dmmu0.page_table\[13\]\[11\] dmmu0.page_table\[14\]\[11\]
+ dmmu0.page_table\[15\]\[11\] _0863_ _0866_ _1221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_40_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5221_ _2332_ _2446_ _2448_ net918 _2467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_59_1990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5152_ _2423_ _0138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6077__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Left_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4103_ _1535_ net272 _1760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3712__I _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5083_ _2140_ _2381_ _2383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4034_ _0813_ _1694_ _1695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5985_ _2782_ _2907_ _2909_ net971 _2911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6621__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4936_ _2294_ _2295_ _1771_ _0050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_25_Left_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_10 net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_21 net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3159__I _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4867_ _2249_ _0027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6001__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input293_I ic0_mem_data[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6606_ _0179_ clknet_leaf_24_core_clock immu_0.page_table\[1\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3818_ _1485_ net665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4798_ _2140_ _2207_ _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3366__A1 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6771__CLK clknet_leaf_99_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6537_ _0110_ clknet_leaf_5_core_clock immu_0.page_table\[7\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3749_ _1405_ _1408_ _1418_ _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6468_ _0041_ clknet_leaf_25_core_clock dmmu0.page_table\[8\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4315__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5419_ _2583_ _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6399_ _0781_ clknet_leaf_0_core_clock immu_0.page_table\[15\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Left_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3669__A2 net375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5291__A1 _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_84_2751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5043__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_2183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_2036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_2047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5594__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5346__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3357__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_2566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3747__I3 _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3109__A1 net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6059__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3532__I _1265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4609__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5806__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_6_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_2016 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6644__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_1102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5770_ _2785_ _0394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5585__A2 _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6794__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4721_ _2162_ _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4652_ _2103_ _2108_ _2110_ immu_1.page_table\[12\]\[9\] _2120_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3348__A1 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3603_ _1302_ net382 _1303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput30 c0_o_mem_data[10] net30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput41 c0_o_mem_data[6] net41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput52 c0_o_mem_high_addr[7] net52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_1531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4583_ _2059_ _2075_ _2077_ net1081 _2080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput63 c0_o_req_addr[13] net63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_1591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput74 c0_o_req_addr[9] net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6322_ _0704_ clknet_leaf_70_core_clock dmmu1.page_table\[14\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_1916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput85 c0_sr_bus_addr[3] net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3534_ _1266_ net553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_57_1927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput96 c0_sr_bus_data_o[1] net96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6253_ _0635_ clknet_leaf_86_core_clock immu_1.page_table\[5\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3465_ _0841_ _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_38_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5204_ _2456_ _0157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6184_ _3023_ _0570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3396_ _0894_ _1128_ _1137_ _1138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3520__A1 net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5135_ _1789_ _2412_ _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4538__I net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input139_I c1_o_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5066_ _2373_ _0102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5273__A1 net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4017_ _1301_ _1678_ _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3823__A2 _1489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input306_I ic0_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5025__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5369__I _2554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5968_ _2900_ _0477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3587__A1 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4784__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4919_ _1994_ _2260_ _2262_ dmmu0.page_table\[8\]\[11\] _2282_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5899_ _2786_ _2856_ _2858_ net923 _2862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3434__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6517__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4839__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3106__A4 net51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput401 inner_wb_i_dat[6] net401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_output525_I net525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6667__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_79_core_clock clknet_4_11__leaf_core_clock clknet_leaf_79_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_67_2223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3814__A2 net705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_63_2109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_2009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5567__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5319__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4527__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6197__CLK clknet_leaf_6_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A3 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3750__A1 _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3750__B2 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3463__S _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3250_ dmmu1.page_table\[1\]\[4\] _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_33_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3181_ _0915_ _0924_ _0929_ _0895_ _0930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__5255__A1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6940_ _0513_ clknet_leaf_59_core_clock dmmu1.page_table\[2\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _0444_ clknet_leaf_55_core_clock dmmu1.page_table\[7\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_46_1606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5007__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5822_ _2047_ _2801_ _2803_ net777 _2816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3569__A1 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5753_ _2773_ _0389_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4704_ _2101_ _2139_ _2142_ net741 _2151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5684_ _2067_ _2726_ _2728_ net1102 _2735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4635_ _2111_ _0742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_66_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _1863_ _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_48_1984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6305_ _0687_ clknet_leaf_89_core_clock immu_1.page_table\[3\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3517_ _0905_ _1254_ _1255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4497_ _1864_ _2014_ _2016_ immu_1.page_table\[3\]\[7\] _2024_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_40_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input256_I dcache_wb_o_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6236_ _0618_ clknet_leaf_83_core_clock immu_1.page_table\[2\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3448_ net154 dmmu1.long_off_reg\[4\] _1188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4297__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6167_ _1535_ net255 _1895_ _3014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3379_ net47 dmmu0.long_off_reg\[2\] _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5118_ _2269_ _2398_ _2400_ immu_0.page_table\[6\]\[3\] _2404_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6098_ _2973_ _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_1668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5246__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5049_ _2328_ _2352_ _2354_ net789 _2363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3352__S0 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5549__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_102_core_clock_I clknet_4_3__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4757__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5827__I _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3548__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4221__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output475_I net475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3980__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3407__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5182__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3791__B _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3732__A1 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5562__I _2665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5485__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_52_core_clock_I clknet_4_13__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput220 dcache_mem_o_data[15] net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3082__I _0843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput231 dcache_wb_adr[0] net231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput242 dcache_wb_adr[1] net242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput253 dcache_wb_adr[8] net253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput264 dcache_wb_o_dat[2] net264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput275 dcache_wb_we net275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput286 ic0_mem_data[18] net286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput297 ic0_mem_data[28] net297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5788__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3799__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3894__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6832__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4420_ _1973_ _1977_ _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_41_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5712__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3723__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4351_ _1861_ _1927_ _1929_ immu_1.page_table\[5\]\[6\] _1936_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3302_ dmmu1.page_table\[8\]\[5\] dmmu1.page_table\[9\]\[5\] dmmu1.page_table\[10\]\[5\]
+ dmmu1.page_table\[11\]\[5\] _0908_ _0910_ _1047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_7070_ net342 net495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_10_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4282_ _1769_ _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XANTENNA__4279__A2 net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6982__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6021_ _2788_ _2924_ _2926_ dmmu1.page_table\[3\]\[4\] _2931_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3233_ dmmu1.page_table\[4\]\[3\] dmmu1.page_table\[5\]\[3\] dmmu1.page_table\[6\]\[3\]
+ dmmu1.page_table\[7\]\[3\] _0899_ _0902_ _0980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_24_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_2044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3164_ _0904_ _0913_ _0895_ _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_59_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5228__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6212__CLK clknet_leaf_97_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3095_ _0840_ _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_72_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _0496_ clknet_leaf_56_core_clock dmmu1.page_table\[3\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__A2 _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6854_ _0427_ clknet_leaf_14_core_clock dmmu0.page_table\[1\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6362__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5805_ _2807_ _0407_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6785_ _0358_ clknet_leaf_52_core_clock dmmu1.page_table\[13\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4203__A2 _1834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3997_ _1440_ _1658_ _1659_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4551__I _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5736_ _2059_ _2760_ _2762_ dmmu1.page_table\[11\]\[2\] _2765_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5951__A2 _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_6_0_core_clock clknet_0_core_clock clknet_3_6_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_72_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3962__A1 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_2059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5667_ _2724_ _0352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input373_I ic1_wb_adr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4618_ _2099_ _0737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5598_ _2453_ _2681_ _2684_ dmmu0.page_table\[6\]\[2\] _2687_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4506__A3 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input67_I c0_o_req_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4911__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4549_ _2057_ _2053_ _2055_ net795 _2058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_2092 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6219_ _0601_ clknet_leaf_90_core_clock immu_1.page_table\[7\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5219__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4690__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7102__I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4978__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6705__CLK clknet_leaf_70_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3876__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output592_I net592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_2058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6855__CLK clknet_leaf_100_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_2115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5155__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3556__I1 net35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4902__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6235__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__CLK clknet_leaf_73_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5630__A1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4433__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3920_ _1375_ _1583_ _1584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_1369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3851_ _1515_ _1516_ _1446_ _1517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5394__B1 _2554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6570_ _0143_ clknet_leaf_7_core_clock immu_0.page_table\[4\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3782_ net705 _1447_ _1450_ _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_27_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5933__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5521_ _2529_ _2630_ _2632_ dmmu0.page_table\[13\]\[9\] _2642_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_82_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_1618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5452_ _2602_ _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_2_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput502 net502 c1_i_req_data[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4044__S1 _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4403_ _1861_ _1957_ _1959_ net945 _1966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput513 net513 c1_i_req_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput524 net524 dcache_mem_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5383_ _2562_ _0230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput535 net535 dcache_mem_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput546 net546 dcache_mem_i_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput557 net557 dcache_mem_i_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7122_ net67 net590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput568 net568 dcache_wb_i_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4334_ _1925_ _0627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput579 net579 dcache_wb_i_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7053_ net290 net441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4265_ _1858_ _1876_ _1878_ immu_1.page_table\[7\]\[5\] _1884_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_10__f_core_clock clknet_3_5_0_core_clock clknet_4_10__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4121__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6004_ _2920_ _0493_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3216_ _0962_ _0963_ _0912_ _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4196_ net187 net186 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6728__CLK clknet_leaf_44_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4672__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3147_ _0896_ _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_input121_I c1_o_mem_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input219_I dcache_mem_o_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3078_ _0819_ _0820_ _0840_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_49_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3858__S1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6906_ _0479_ clknet_leaf_59_core_clock dmmu1.page_table\[5\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_2069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6837_ _0410_ clknet_leaf_51_core_clock dmmu1.page_table\[9\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3098__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6768_ _0341_ clknet_leaf_41_core_clock dmmu0.page_table\[5\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3935__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5719_ _2754_ _0374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6699_ _0272_ clknet_leaf_34_core_clock dmmu0.page_table\[4\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5688__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3538__I1 net41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6258__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold260 dmmu0.page_table\[4\]\[2\] net994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3163__A2 _0911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold271 dmmu0.page_table\[11\]\[9\] net1005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold282 dmmu0.page_table\[14\]\[6\] net1016 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold293 dmmu0.page_table\[10\]\[6\] net1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_79_1516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output438_I net438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6101__A2 _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5860__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_1858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4415__A2 _1972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5612__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__I1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3849__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5376__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5128__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3963__C _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4026__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3529__I1 net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4351__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4103__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4050_ net10 immu_0.high_addr_off\[5\] _1710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 c0_o_instr_long_addr[1] net6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_1909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4952_ _2271_ _2299_ _2302_ dmmu0.page_table\[7\]\[4\] _2307_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_52_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3903_ _1463_ immu_0.page_table\[11\]\[5\] _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4883_ _2257_ _0035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6159__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3834_ _1499_ _1500_ _1439_ _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6622_ _0195_ clknet_leaf_20_core_clock immu_0.page_table\[0\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6553_ _0126_ clknet_leaf_27_core_clock immu_0.page_table\[6\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3765_ _1416_ _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_67_1420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5504_ _2633_ _0280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_82_1918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6484_ _0057_ clknet_leaf_16_core_clock dmmu0.page_table\[7\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3696_ net314 _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_28_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5435_ _2592_ _0252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3145__A2 net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input169_I c1_o_req_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ _1781_ _1977_ _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_61_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6550__CLK clknet_leaf_6_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4893__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7105_ net396 net573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4317_ _1849_ _1911_ _1914_ net934 _1917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5297_ net103 _2502_ _2504_ immu_0.page_table\[0\]\[8\] _2512_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_10_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6095__A1 net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7036_ net303 net454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input336_I ic1_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4248_ net190 _1872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__5842__A1 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4179_ net103 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_39_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_2690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5358__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_14_Right_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_1586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3556__S _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3783__C _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4581__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4008__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_2494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4333__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3767__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_2369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_23_Right_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4636__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3090__I _0847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5061__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3072__A1 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Right_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6423__CLK clknet_leaf_112_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3550_ net137 net32 _1267_ _1275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6573__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_2002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3481_ dmmu0.page_table\[8\]\[11\] dmmu0.page_table\[9\]\[11\] dmmu0.page_table\[10\]\[11\]
+ dmmu0.page_table\[11\]\[11\] _0871_ _0867_ _1220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_45_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5220_ _2466_ _0163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_59_1980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_59_1991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_41_Right_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5521__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_2068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1946 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5151_ _2275_ _2414_ _2416_ net900 _2423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_55_1877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6077__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4102_ _1350_ net326 _1360_ _1759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5082_ _2381_ _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_36_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5824__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4033_ _1502_ _1688_ _1693_ net705 _1694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_75_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__I _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3868__C _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_50_Right_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5984_ _2910_ _0483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4935_ _1796_ _2290_ _2291_ _1845_ _2295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_11 net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_22 net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4866_ _1806_ _2242_ _2244_ dmmu0.page_table\[9\]\[4\] _2249_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_1526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6001__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6916__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_107_core_clock_I clknet_4_2__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6605_ _0178_ clknet_leaf_18_core_clock immu_0.page_table\[1\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3817_ net236 _1484_ _1360_ _1485_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4797_ _2207_ _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_55_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input286_I ic0_mem_data[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3748_ _1408_ _1417_ _1418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6536_ _0109_ clknet_leaf_10_core_clock immu_0.page_table\[8\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6467_ _0040_ clknet_leaf_31_core_clock dmmu0.page_table\[8\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3679_ _1348_ net377 _1353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4315__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5418_ _2300_ _2581_ _2583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6398_ _0780_ clknet_leaf_0_core_clock immu_0.page_table\[15\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4866__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5349_ _2543_ _0215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_69_core_clock clknet_4_12__leaf_core_clock clknet_leaf_69_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5666__I1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_57_core_clock_I clknet_4_14__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5291__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3921__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6446__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3778__C _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5579__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7110__I net401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_2627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5043__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_2173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_2037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_2048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_2059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_2545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_2556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3109__A2 _0858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6059__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5806__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4609__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5282__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3293__A1 _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3045__A1 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_48_1670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4720_ _1800_ _2157_ _2159_ immu_0.page_table\[15\]\[2\] _2162_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_29_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4651_ _2119_ _0750_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3602_ _1301_ _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput20 c0_o_mem_addr[1] net20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput31 c0_o_mem_data[11] net31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5742__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3979__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4582_ _2079_ _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput42 c0_o_mem_data[7] net42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput53 c0_o_mem_long_mode net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput64 c0_o_req_addr[14] net64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3533_ net144 net39 _0850_ _1266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput75 c0_o_req_ppl_submit net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6321_ _0703_ clknet_leaf_98_core_clock dmmu1.page_table\[14\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput86 c0_sr_bus_addr[4] net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_1917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput97 c0_sr_bus_data_o[2] net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_1939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6252_ _0634_ clknet_leaf_89_core_clock immu_1.page_table\[5\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3464_ _1203_ net531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5203_ _2455_ _2447_ _2449_ immu_0.page_table\[3\]\[3\] _2456_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6183_ dmmu1.long_off_reg\[6\] _1861_ _3016_ _3023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3395_ _0915_ _1131_ _1136_ _0894_ _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5134_ _2205_ _2296_ _2412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_77_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6469__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5065_ _2269_ _2367_ _2369_ net922 _2373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4016_ _1378_ _1672_ _1677_ _1381_ _1678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__5273__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3284__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4554__I _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input201_I c1_sr_bus_data_o[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5025__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3036__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5967_ _2794_ _2890_ _2892_ net792 _2900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4784__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3587__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4918_ _2281_ _0046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_1293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5898_ _2861_ _0446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input97_I c0_sr_bus_data_o[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4849_ _1994_ _2223_ _2225_ dmmu0.page_table\[10\]\[11\] _2238_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4536__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6519_ _0092_ clknet_leaf_4_core_clock immu_0.page_table\[9\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_2420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3834__S _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4839__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7105__I net396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput402 inner_wb_i_dat[7] net402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_67_2224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3275__A1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4527__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3750__A2 _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3543__I _1271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3180_ _0926_ _0928_ _0915_ _0929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5255__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_53_Left_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3266__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4463__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6870_ _0443_ clknet_leaf_68_core_clock dmmu1.page_table\[8\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_46_1607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5007__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5821_ _2815_ _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3569__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5963__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ _2105_ _2759_ _2761_ net855 _2773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4703_ _2150_ _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5683_ _2734_ _0358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_62_Left_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4634_ _2051_ _2108_ _2110_ net825 _2111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4565_ _2068_ _0715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3881__C _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6304_ _0686_ clknet_leaf_82_core_clock immu_1.page_table\[3\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3516_ dmmu1.page_table\[8\]\[12\] dmmu1.page_table\[9\]\[12\] dmmu1.page_table\[10\]\[12\]
+ dmmu1.page_table\[11\]\[12\] _0886_ net121 _1254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_12_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4496_ _2023_ _0691_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Right_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6291__CLK clknet_leaf_101_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6235_ _0617_ clknet_leaf_80_core_clock immu_1.page_table\[2\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3447_ net155 dmmu1.long_off_reg\[5\] _1187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input151_I c1_o_mem_high_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input249_I dcache_wb_adr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3378_ net47 dmmu0.long_off_reg\[2\] _1120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6166_ _3013_ _0562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_71_Left_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5117_ _2403_ _0123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6097_ net200 _2957_ _2959_ net835 _2973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5246__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5048_ _2362_ _0095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3257__A1 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input12_I c0_o_instr_long_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3352__S1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6999_ _0572_ clknet_leaf_106_core_clock icore_sregs.c1_disable vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4757__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Left_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4509__A1 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5706__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5182__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_2016 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6634__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3732__A2 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output635_I net635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5485__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput210 c1_sr_bus_we net210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3496__A1 net51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6784__CLK clknet_leaf_46_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput221 dcache_mem_o_data[1] net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput232 dcache_wb_adr[10] net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput243 dcache_wb_adr[20] net243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput254 dcache_wb_adr[9] net254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput265 dcache_wb_o_dat[3] net265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput276 ic0_mem_ack net276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_1709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput287 ic0_mem_data[19] net287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput298 ic0_mem_data[29] net298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3248__A1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3799__A2 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4350_ _1935_ _0633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_50_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3301_ _0907_ _1045_ _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4281_ _1893_ _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_26_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6020_ _2930_ _0499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3232_ _0977_ _0978_ _0884_ _0979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__3487__A1 _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_2034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input4_I c0_o_icache_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3163_ _0907_ _0911_ _0912_ _0913_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_55_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5228__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3094_ _0849_ net537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3222__B _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6922_ _0495_ clknet_leaf_64_core_clock dmmu1.page_table\[4\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6507__CLK clknet_leaf_2_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6853_ _0426_ clknet_leaf_43_core_clock dmmu0.page_table\[1\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5804_ _2784_ _2802_ _2804_ dmmu1.page_table\[9\]\[2\] _2807_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6784_ _0357_ clknet_leaf_46_core_clock dmmu1.page_table\[13\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3996_ immu_1.page_table\[8\]\[8\] immu_1.page_table\[9\]\[8\] immu_1.page_table\[10\]\[8\]
+ immu_1.page_table\[11\]\[8\] _1441_ _1540_ _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_50_1864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5735_ _2764_ _0380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6657__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input199_I c1_sr_bus_data_o[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5666_ dmmu0.long_off_reg\[7\] _1815_ _2716_ _2724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5164__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4617_ _2067_ _2090_ _2092_ immu_1.page_table\[13\]\[6\] _2099_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5597_ _2686_ _0320_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input366_I ic1_wb_adr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4911__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4548_ _1845_ _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_13_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6113__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3183__I net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4479_ _1838_ _1874_ _1891_ _2013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6218_ _0600_ clknet_leaf_90_core_clock immu_1.page_table\[7\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3478__A1 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6149_ _1848_ _3000_ _3002_ net1073 _3005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5219__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4427__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4978__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3650__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4742__I _2174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5927__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_2015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output585_I net585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3402__A1 net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5155__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__I _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3308__I2 dmmu0.page_table\[14\]\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3469__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4666__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2016 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_2084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5091__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3641__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3850_ immu_1.page_table\[4\]\[4\] immu_1.page_table\[5\]\[4\] immu_1.page_table\[6\]\[4\]
+ immu_1.page_table\[7\]\[4\] _1441_ _1442_ _1516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_15_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1072 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3781_ _1440_ _1448_ _1449_ _1444_ _1415_ _1450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__5394__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3268__I net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5520_ _2641_ _0288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5451_ _1834_ _2601_ _2602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_1960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_2033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_2093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4402_ _1965_ _0655_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput503 net503 c1_i_req_data[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput514 net514 c1_i_req_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput525 net525 dcache_mem_addr[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5382_ _2461_ _2553_ _2555_ dmmu0.page_table\[11\]\[6\] _2562_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput536 net536 dcache_mem_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput547 net547 dcache_mem_i_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7121_ net66 net589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput558 net558 dcache_mem_i_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4333_ _1870_ _1910_ _1913_ immu_1.page_table\[2\]\[10\] _1925_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput569 net569 dcache_wb_i_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5449__A2 _1836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4264_ _1883_ _0599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7052_ net289 net440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3215_ dmmu1.page_table\[8\]\[2\] dmmu1.page_table\[9\]\[2\] dmmu1.page_table\[10\]\[2\]
+ dmmu1.page_table\[11\]\[2\] _0899_ _0902_ _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6003_ _2851_ _2906_ _2908_ dmmu1.page_table\[4\]\[10\] _2920_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4121__A2 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4195_ net195 _1830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3146_ net122 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4409__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3880__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3077_ _0839_ net473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_2015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input114_I c1_o_instr_long_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6905_ _0478_ clknet_leaf_61_core_clock dmmu1.page_table\[5\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6836_ _0409_ clknet_leaf_52_core_clock dmmu1.page_table\[9\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5909__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6767_ _0340_ clknet_leaf_49_core_clock dmmu0.page_table\[5\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3979_ immu_0.page_table\[8\]\[7\] immu_0.page_table\[9\]\[7\] immu_0.page_table\[10\]\[7\]
+ immu_0.page_table\[11\]\[7\] _1487_ _1390_ _1642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_50_1683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5718_ _2101_ _2743_ _2745_ net815 _2754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6698_ _0271_ clknet_leaf_36_core_clock dmmu0.page_table\[4\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5137__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5649_ _2714_ _0344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5688__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4896__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold250 immu_0.page_table\[12\]\[9\] net984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold261 immu_0.page_table\[12\]\[0\] net995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold272 dmmu1.page_table\[1\]\[1\] net1006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold283 dmmu0.page_table\[9\]\[0\] net1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold294 immu_0.page_table\[11\]\[2\] net1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_79_1528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4648__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7113__I net404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5860__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3871__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output500_I net500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6822__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5073__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5612__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3623__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5376__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6972__CLK clknet_leaf_64_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3088__I _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3226__I1 _0972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3482__S0 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_64_core_clock_I clknet_4_11__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5128__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6202__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3234__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4351__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4103__A2 net272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3551__I _1275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput7 c0_o_instr_long_addr[2] net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4951_ _2306_ _0054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_52_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3902_ _1385_ immu_0.page_table\[10\]\[5\] _1567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4882_ _1996_ _2241_ _2243_ dmmu0.page_table\[9\]\[12\] _2257_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_51_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6621_ _0194_ clknet_leaf_16_core_clock immu_0.page_table\[0\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3833_ immu_1.page_table\[0\]\[3\] immu_1.page_table\[1\]\[3\] immu_1.page_table\[2\]\[3\]
+ immu_1.page_table\[3\]\[3\] _1435_ _1469_ _1500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_55_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6552_ _0125_ clknet_leaf_21_core_clock immu_0.page_table\[6\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3764_ _1410_ _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_27_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3473__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5503_ _2444_ _2630_ _2632_ net1072 _2633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6483_ _0056_ clknet_leaf_32_core_clock dmmu0.page_table\[7\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3726__I _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3695_ _1363_ _1364_ _1365_ net662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_14_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5434_ _2463_ _2582_ _2584_ net940 _2592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3225__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4878__B1 _2243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5365_ _2551_ _0223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7104_ net389 net566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_1687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4316_ _1916_ _0618_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5296_ _2511_ _0194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6095__A2 _2957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4557__I _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7035_ net302 net453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_59_core_clock clknet_4_15__leaf_core_clock clknet_leaf_59_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4247_ _1871_ _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6845__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input231_I dcache_wb_adr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input329_I ic0_wb_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5842__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4178_ _1816_ _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_1403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3129_ _0878_ _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6995__CLK clknet_leaf_97_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4802__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_2680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_2691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6819_ _0392_ clknet_leaf_50_core_clock dmmu1.page_table\[10\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5358__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6225__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4581__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7108__I net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_98_core_clock clknet_4_9__leaf_core_clock clknet_leaf_98_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_76_2484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6375__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_2495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_2004 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3767__S1 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4097__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3844__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_2092 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3072__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4021__A1 net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6718__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_1774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3480_ _0841_ _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_1914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5521__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6868__CLK clknet_leaf_67_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5150_ _2422_ _0137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_55_1867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6077__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4101_ _1348_ net380 _1758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_1379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5081_ _1790_ _2297_ _2381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_36_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4088__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5285__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4032_ _1415_ _1690_ _1692_ _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_79_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5037__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5983_ _2776_ _2907_ _2909_ net944 _2910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6248__CLK clknet_leaf_90_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4934_ net407 _2293_ _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4045__C _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4865_ _2248_ _0026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_12 net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_23 net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6001__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6604_ _0177_ clknet_leaf_7_core_clock immu_0.page_table\[1\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3816_ _1422_ _1459_ _1468_ _1473_ _1483_ _1484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__4012__A1 _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6398__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ _1790_ _2206_ _2207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_43_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6535_ _0108_ clknet_leaf_5_core_clock immu_0.page_table\[8\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3747_ _1411_ _1412_ _1413_ _1414_ _1415_ _1416_ _1417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_42_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input181_I c1_sr_bus_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input279_I ic0_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6466_ _0039_ clknet_leaf_32_core_clock dmmu0.page_table\[8\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3678_ _1349_ _1351_ _1352_ net681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4315__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5417_ _2581_ _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6397_ _0779_ clknet_leaf_112_core_clock immu_0.page_table\[15\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5348_ _2457_ _2536_ _2538_ net867 _2543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input42_I c0_o_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3191__I _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4079__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5279_ _2501_ _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_39_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3826__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_2731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3921__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_2742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5579__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_80_2617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4251__A1 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_2049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output498_I net498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5200__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_2546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5503__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6059__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5267__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5806__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5019__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_48_1660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3045__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__CLK clknet_leaf_26_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4650_ _2101_ _2108_ _2110_ net983 _2119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_56_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3601_ icache_arbiter.o_sel_sig _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
Xinput10 c0_o_instr_long_addr[5] net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5742__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput21 c0_o_mem_addr[2] net21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput32 c0_o_mem_data[12] net32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_24_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3979__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4581_ _2057_ _2075_ _2077_ immu_1.page_table\[14\]\[1\] _2079_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput43 c0_o_mem_data[8] net43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6690__CLK clknet_leaf_92_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput54 c0_o_mem_req net54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6320_ _0702_ clknet_leaf_71_core_clock dmmu1.page_table\[14\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3532_ _1265_ net552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput65 c0_o_req_addr[15] net65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput76 c0_sr_bus_addr[0] net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_3_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput87 c0_sr_bus_addr[5] net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput98 c0_sr_bus_data_o[3] net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_57_1929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6251_ _0633_ clknet_leaf_87_core_clock immu_1.page_table\[5\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3463_ _1186_ _1202_ _0884_ _1203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5202_ _1802_ _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6182_ _3022_ _0569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3394_ net123 _1133_ _1135_ _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_62_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5133_ _2411_ _0131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_4_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5064_ _2372_ _0101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3808__A1 _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4015_ _1377_ _1674_ _1676_ _1677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_79_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4481__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5966_ _2899_ _0476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3036__A2 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5430__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_106_core_clock clknet_4_2__leaf_core_clock clknet_leaf_106_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4917_ _1821_ _2260_ _2262_ net1048 _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4784__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5981__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ _2784_ _2856_ _2858_ net989 _2861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input396_I inner_wb_i_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4848_ _2237_ _0020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3419__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4779_ _2197_ _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6518_ _0091_ clknet_leaf_9_core_clock immu_0.page_table\[9\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_73_2410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_1508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ _0022_ clknet_leaf_102_core_clock dmmu0.page_table\[10\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_1688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3135__B _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput403 inner_wb_i_dat[8] net403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6413__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_2214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_2236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7121__I net66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_2002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3822__I1 _1488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4527__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5724__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_33_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6906__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4463__A1 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7031__I net406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3266__A2 _0994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_1608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5820_ _2105_ _2801_ _2803_ net1045 _2815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5751_ _2772_ _0388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5963__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _2069_ _2139_ _2142_ net962 _2150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5682_ _2065_ _2726_ _2728_ net865 _2734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4633_ _2109_ _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_72_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4074__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4564_ _2067_ _2053_ _2055_ net987 _2068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_83_1855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3821__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6303_ _0685_ clknet_leaf_83_core_clock immu_1.page_table\[3\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3515_ _1251_ _1252_ _0896_ _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_1385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4495_ _1861_ _2014_ _2016_ net775 _2023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3734__I net366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5479__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6234_ _0616_ clknet_leaf_96_core_clock immu_1.page_table\[0\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3446_ _1179_ _1185_ _1186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6165_ _2851_ _2999_ _3001_ immu_1.page_table\[8\]\[10\] _3013_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3377_ net53 _0859_ _1119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_input144_I c1_o_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5116_ _2267_ _2398_ _2400_ immu_0.page_table\[6\]\[2\] _2403_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6586__CLK clknet_leaf_24_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6096_ _2972_ _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5047_ _2277_ _2352_ _2354_ immu_0.page_table\[9\]\[7\] _2362_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input311_I ic0_wb_adr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1946 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6998_ _0571_ clknet_leaf_98_core_clock dmmu1.long_off_reg\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4757__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5949_ _1828_ _1873_ _2030_ _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_48_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4509__A2 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5706__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5182__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_69_core_clock_I clknet_4_12__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7116__I net392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6131__A1 net559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6929__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output628_I net628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput200 c1_sr_bus_data_o[12] net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput211 core_reset net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xinput222 dcache_mem_o_data[2] net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput233 dcache_wb_adr[11] net233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput244 dcache_wb_adr[21] net244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput255 dcache_wb_cyc net255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput266 dcache_wb_o_dat[4] net266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput277 ic0_mem_data[0] net277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput288 ic0_mem_data[1] net288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput299 ic0_mem_data[2] net299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4445__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5642__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6309__CLK clknet_leaf_96_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4056__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6459__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3982__C _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3803__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3184__A1 net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4381__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3300_ dmmu1.page_table\[12\]\[5\] dmmu1.page_table\[13\]\[5\] dmmu1.page_table\[14\]\[5\]
+ dmmu1.page_table\[15\]\[5\] _0888_ _0910_ _1045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_22_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4280_ _1838_ _1891_ _1892_ _1893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_26_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3231_ _0879_ _0883_ _0978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_1260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_2046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3162_ net123 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_20_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3093_ net129 net24 _0842_ _0849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_71_core_clock_I clknet_4_9__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6921_ _0494_ clknet_leaf_65_core_clock dmmu1.page_table\[4\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6189__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6852_ _0425_ clknet_leaf_37_core_clock dmmu0.page_table\[1\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5803_ _2806_ _0406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6783_ _0356_ clknet_leaf_48_core_clock dmmu1.page_table\[13\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4739__A2 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3995_ _1655_ _1656_ _1439_ _1657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5734_ _2057_ _2760_ _2762_ net875 _2764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_1985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5665_ _2723_ _0351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_1685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4616_ _2098_ _0736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5164__A2 _2429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5596_ _2451_ _2681_ _2684_ dmmu0.page_table\[6\]\[1\] _2686_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_1750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4547_ _2056_ _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4911__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3464__I _1203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input261_I dcache_wb_o_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input359_I ic1_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6113__A1 _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4478_ _2012_ _0684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6217_ _0599_ clknet_leaf_84_core_clock immu_1.page_table\[7\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3429_ _1154_ _1169_ _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_42_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5872__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6148_ _3004_ _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6079_ _2786_ _2958_ _2960_ net1082 _2964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4427__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5624__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4978__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3650__A2 net242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5927__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6601__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output480_I net480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5155__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6751__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3307__C _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_15__f_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4418__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_2074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5091__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3641__A2 net262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3549__I _1274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6281__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5394__A2 _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3780_ immu_1.page_table\[10\]\[1\] immu_1.page_table\[11\]\[1\] _1404_ _1449_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5450_ _1891_ _1892_ _2599_ _2600_ _2601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_67_1658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4401_ _1858_ _1957_ _1959_ net967 _1965_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput504 net504 c1_i_req_data[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5381_ _2561_ _0229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput515 net515 c1_i_req_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput526 net526 dcache_mem_addr[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput537 net537 dcache_mem_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7120_ net59 net582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput548 net548 dcache_mem_i_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4332_ _1924_ _0626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput559 net559 dcache_mem_req vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_61_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7051_ net287 net438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_49_core_clock clknet_4_13__leaf_core_clock clknet_leaf_49_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4263_ _1855_ _1876_ _1878_ immu_1.page_table\[7\]\[4\] _1883_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__B1 _2820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6002_ _2919_ _0492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3214_ dmmu1.page_table\[0\]\[2\] dmmu1.page_table\[1\]\[2\] dmmu1.page_table\[2\]\[2\]
+ dmmu1.page_table\[3\]\[2\] _0899_ _0931_ _0962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__4121__A3 _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4194_ _1826_ _1828_ _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3145_ net106 net158 _0894_ _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__4409__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5004__I _2336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_2010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5606__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3076_ net220 _0831_ _0839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_1440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6624__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6904_ _0477_ clknet_leaf_61_core_clock dmmu1.page_table\[5\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input107_I c1_o_c_instr_long vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6835_ _0408_ clknet_leaf_49_core_clock dmmu1.page_table\[9\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_1894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5909__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6031__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6766_ _0339_ clknet_leaf_35_core_clock dmmu0.page_table\[5\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3978_ _1375_ _1640_ _1641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3396__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4593__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5717_ _2753_ _0373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6697_ _0270_ clknet_leaf_49_core_clock dmmu0.page_table\[4\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5648_ net95 _2698_ _2700_ net985 _2714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_88_core_clock clknet_4_10__leaf_core_clock clknet_leaf_88_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6185__I1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input72_I c0_o_req_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ _2101_ _2664_ _2666_ net808 _2675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4896__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold240 dmmu1.page_table\[15\]\[11\] net974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold251 dmmu0.page_table\[5\]\[12\] net985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold262 dmmu0.page_table\[5\]\[8\] net996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold273 dmmu0.page_table\[10\]\[5\] net1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold284 dmmu1.page_table\[2\]\[3\] net1018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold295 dmmu0.page_table\[6\]\[7\] net1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4648__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5073__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3623__A2 net268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4820__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5376__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3482__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5128__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3234__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5836__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3311__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6647__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 c0_o_instr_long_addr[3] net8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_1938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4950_ _2269_ _2299_ _2302_ dmmu0.page_table\[7\]\[3\] _2306_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_1613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6797__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3901_ _1564_ _1565_ _1367_ _1566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4881_ _2256_ _0034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6013__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6620_ _0193_ clknet_leaf_19_core_clock immu_0.page_table\[0\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3832_ immu_1.page_table\[4\]\[3\] immu_1.page_table\[5\]\[3\] immu_1.page_table\[6\]\[3\]
+ immu_1.page_table\[7\]\[3\] _1435_ _1469_ _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_6_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3378__A1 net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6551_ _0124_ clknet_leaf_26_core_clock immu_0.page_table\[6\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3763_ _1375_ _1428_ _1431_ _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_15_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5502_ _2631_ _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3473__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_2009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6482_ _0055_ clknet_leaf_32_core_clock dmmu0.page_table\[7\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3694_ _1337_ net233 _1365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_1417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4327__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5433_ _2591_ _0251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3225__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4878__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5364_ _1996_ _2535_ _2537_ net861 _2551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_80_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7103_ net211 net563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4315_ _1846_ _1911_ _1914_ immu_1.page_table\[2\]\[1\] _1916_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5295_ _1814_ _2502_ _2504_ immu_0.page_table\[0\]\[7\] _2511_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7034_ net299 net450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4246_ _1870_ _1840_ _1842_ immu_1.page_table\[9\]\[10\] _1871_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4177_ _1815_ _1792_ _1794_ immu_0.page_table\[11\]\[7\] _1816_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input224_I dcache_mem_o_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3128_ net18 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5669__I _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3059_ net227 _0822_ _0830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4802__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3161__S0 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_2670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_2681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3189__I _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _0391_ clknet_leaf_68_core_clock dmmu1.page_table\[11\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5358__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6749_ _0322_ clknet_leaf_35_core_clock dmmu0.page_table\[6\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_2485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_2496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output443_I net443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7124__I net69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5818__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4097__A2 net383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3844__A2 net705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3099__I _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5521__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7034__I net299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_55_1879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4100_ _1755_ _1756_ _1757_ net704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5080_ _2380_ _0109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_10_core_clock_I clknet_4_3__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5285__A1 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4031_ _1416_ _1691_ _1692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_13 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5037__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5982_ _2908_ _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_75_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3599__A1 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4933_ _1796_ _2285_ _2287_ _1845_ _2293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4864_ _1803_ _2242_ _2244_ net914 _2248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_13 net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3815_ _0813_ _1482_ _1483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_24 net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6603_ _0176_ clknet_leaf_19_core_clock immu_0.page_table\[1\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4795_ _2154_ _2205_ _2206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_16_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6534_ _0107_ clknet_leaf_5_core_clock immu_0.page_table\[8\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ net368 _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_43_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6465_ _0038_ clknet_leaf_31_core_clock dmmu0.page_table\[8\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3677_ _1337_ net252 _1352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6812__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input174_I c1_o_req_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5416_ _1977_ _2468_ _2581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6396_ _0778_ clknet_leaf_108_core_clock immu_0.page_table\[15\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5347_ _2542_ _0214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4720__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_2360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input341_I ic1_mem_data[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5278_ _1789_ _1973_ _2501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6962__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input35_I c0_o_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4229_ _1858_ _1841_ _1843_ net936 _1859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_2732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5579__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_2175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4251__A2 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6342__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_inner_730 c1_i_core_int_sreg[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_85_2042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7119__I net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5200__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_2558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3762__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6492__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_1_core_clock_I clknet_4_0__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5267__A1 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3373__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5019__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_76_core_clock_I clknet_4_11__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4778__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4941__I _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1004 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_1649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3557__I _1278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6835__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3600_ _1300_ net427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 c0_o_instr_long_addr[6] net11 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_1750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput22 c0_o_mem_addr[3] net22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4580_ _2078_ _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5742__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput33 c0_o_mem_data[13] net33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_80_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput44 c0_o_mem_data[9] net44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput55 c0_o_mem_sel[0] net55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3531_ net143 net38 _0850_ _1265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4950__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput66 c0_o_req_addr[1] net66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput77 c0_sr_bus_addr[10] net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_1919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput88 c0_sr_bus_addr[6] net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6250_ _0632_ clknet_leaf_85_core_clock immu_1.page_table\[5\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput99 c0_sr_bus_data_o[4] net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3462_ _0894_ _1191_ _1192_ _0895_ _1201_ _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_0_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6985__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3505__A1 _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5201_ _2454_ _0156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4702__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6181_ dmmu1.long_off_reg\[5\] _1858_ _3016_ _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3393_ _0906_ _1134_ _1135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5132_ _2332_ _2397_ _2399_ net818 _2411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6215__CLK clknet_leaf_90_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5063_ _2267_ _2367_ _2369_ net753 _2372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4014_ _1366_ _1675_ _1676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_7__f_core_clock clknet_3_3_0_core_clock clknet_4_7__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_75_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3241__B _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6365__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5965_ _2792_ _2890_ _2892_ dmmu1.page_table\[5\]\[6\] _2899_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3036__A3 _0815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5430__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_1885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4916_ _2280_ _0045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5896_ _2860_ _0445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5981__A2 _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4847_ _1821_ _2223_ _2225_ dmmu0.page_table\[10\]\[10\] _2237_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3419__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input291_I ic0_mem_data[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input389_I inner_wb_i_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5194__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4778_ _1803_ _2191_ _2193_ immu_0.page_table\[12\]\[3\] _2197_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3729_ _1394_ _1395_ _1398_ _1372_ _1366_ _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_6517_ _0090_ clknet_leaf_7_core_clock immu_0.page_table\[9\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_2400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_2070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6448_ _0021_ clknet_leaf_12_core_clock dmmu0.page_table\[10\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5497__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6379_ _0761_ clknet_leaf_77_core_clock immu_1.page_table\[11\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput404 inner_wb_i_dat[9] net404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_41_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_1318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_67_2215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6708__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_2226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output406_I net406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6858__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3983__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6238__CLK clknet_leaf_91_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6388__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3346__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4999__B1 _2318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4463__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3266__A3 _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5750_ _2103_ _2760_ _2762_ dmmu1.page_table\[11\]\[9\] _2772_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5963__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4701_ _2149_ _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5681_ _2733_ _0357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4632_ _1912_ _2107_ _2109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5176__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4074__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4563_ _1860_ _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_8_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3821__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6302_ _0684_ clknet_leaf_96_core_clock immu_1.page_table\[1\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3514_ dmmu1.page_table\[4\]\[12\] dmmu1.page_table\[5\]\[12\] dmmu1.page_table\[6\]\[12\]
+ dmmu1.page_table\[7\]\[12\] _0886_ _0900_ _1252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4494_ _2022_ _0690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_83_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5479__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6233_ _0615_ clknet_leaf_83_core_clock immu_1.page_table\[0\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3445_ _1180_ _1183_ _1184_ _1185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6164_ _3012_ _0561_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3376_ _0879_ _1112_ _1117_ _0860_ _1118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_5115_ _2402_ _0122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6095_ net199 _2957_ _2959_ net796 _2972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input137_I c1_o_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5046_ _2361_ _0094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input304_I ic0_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6997_ _0570_ clknet_leaf_98_core_clock dmmu1.long_off_reg\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5948_ _2888_ _0469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3965__A1 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5879_ net209 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_29_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4509__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5706__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_1497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4142__A1 net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput201 c1_sr_bus_data_o[1] net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput212 dcache_mem_ack net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_output523_I net523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput223 dcache_mem_o_data[3] net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput234 dcache_wb_adr[12] net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput245 dcache_wb_adr[22] net245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7132__I net62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput256 dcache_wb_o_dat[0] net256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput267 dcache_wb_o_dat[5] net267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3328__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput278 ic0_mem_data[10] net278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput289 ic0_mem_data[20] net289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4445__A2 _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5642__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6680__CLK clknet_leaf_40_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Left_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3500__S0 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4056__S1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4905__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3835__I _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3803__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4381__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_39_core_clock clknet_4_6__leaf_core_clock clknet_leaf_39_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3230_ _0975_ _0976_ _0938_ _0977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3161_ dmmu1.page_table\[0\]\[0\] dmmu1.page_table\[1\]\[0\] dmmu1.page_table\[2\]\[0\]
+ dmmu1.page_table\[3\]\[0\] _0908_ _0910_ _0911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__7042__I net278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3092_ _0848_ net536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6920_ _0493_ clknet_leaf_65_core_clock dmmu1.page_table\[4\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6851_ _0424_ clknet_leaf_41_core_clock dmmu0.page_table\[1\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5802_ _2782_ _2802_ _2804_ net889 _2806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3994_ immu_1.page_table\[0\]\[8\] immu_1.page_table\[1\]\[8\] immu_1.page_table\[2\]\[8\]
+ immu_1.page_table\[3\]\[8\] _1404_ _1540_ _1656_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6782_ _0355_ clknet_leaf_48_core_clock dmmu1.page_table\[13\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3947__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5733_ _2763_ _0379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5149__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5664_ dmmu0.long_off_reg\[6\] _1812_ _2716_ _2723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_78_core_clock clknet_4_11__leaf_core_clock clknet_leaf_78_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_44_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4615_ _2065_ _2090_ _2092_ immu_1.page_table\[13\]\[5\] _2098_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5595_ _2685_ _0319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3745__I net369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4546_ _2051_ _2053_ _2055_ net869 _2056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_83_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6553__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4477_ net198 _1998_ _2000_ immu_1.page_table\[1\]\[10\] _2012_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6113__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input254_I dcache_wb_adr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4124__A1 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5321__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6216_ _0598_ clknet_leaf_91_core_clock immu_1.page_table\[7\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3428_ _1159_ _1168_ _0821_ _1169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5872__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_1383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6147_ _1845_ _3000_ _3002_ net954 _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3480__I _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3359_ _0938_ _1101_ _0958_ _1102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6078_ _2963_ _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5624__A1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4427__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5029_ _1790_ _2240_ _2351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_68_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5388__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5927__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_2017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7127__I net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4363__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output640_I net640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4666__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_15_core_clock_I clknet_4_6__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5091__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6426__CLK clknet_leaf_110_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3929__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6576__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7037__I net304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4400_ _1964_ _0654_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_84_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5551__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3788__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5380_ _2459_ _2553_ _2555_ dmmu0.page_table\[11\]\[5\] _2561_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_84_1973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput505 net505 c1_i_req_data[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput516 net516 c1_i_req_data_valid vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_50_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput527 net527 dcache_mem_addr[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4331_ _1868_ _1911_ _1914_ immu_1.page_table\[2\]\[9\] _1924_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput538 net538 dcache_mem_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput549 net549 dcache_mem_i_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5780__I _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7050_ net286 net437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4106__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4262_ _1882_ _0598_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5854__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6001_ _2849_ _2907_ _2909_ net951 _2919_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3213_ _0959_ _0960_ _0884_ _0961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_43_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4193_ _1827_ net181 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_78_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3144_ net158 _0893_ _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__3960__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4409__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5606__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5457__I1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3075_ _0838_ net472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6903_ _0476_ clknet_leaf_56_core_clock dmmu1.page_table\[5\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Left_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6834_ _0407_ clknet_leaf_49_core_clock dmmu1.page_table\[9\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5909__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6031__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6765_ _0338_ clknet_leaf_14_core_clock dmmu0.page_table\[5\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3977_ immu_0.page_table\[12\]\[7\] immu_0.page_table\[13\]\[7\] immu_0.page_table\[14\]\[7\]
+ immu_0.page_table\[15\]\[7\] _1487_ _1390_ _1640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4593__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3396__A2 _1128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5716_ _2069_ _2743_ _2745_ net862 _2753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6696_ _0269_ clknet_leaf_34_core_clock dmmu0.page_table\[4\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5647_ _2713_ _0343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input371_I ic1_wb_adr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4345__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3779__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5578_ _2674_ _0313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input65_I c0_o_req_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold230 dmmu0.page_table\[1\]\[10\] net964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4896__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Left_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold241 immu_1.page_table\[2\]\[7\] net975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4529_ _1866_ _2033_ _2035_ dmmu1.page_table\[14\]\[8\] _2044_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold252 dmmu1.page_table\[10\]\[8\] net986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold263 dmmu0.page_table\[13\]\[5\] net997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold274 immu_1.page_table\[5\]\[5\] net1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold285 immu_0.page_table\[13\]\[10\] net1019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold296 dmmu1.page_table\[7\]\[1\] net1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4648__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_6_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7179_ net398 net651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_6_core_clock_I clknet_4_1__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3871__A3 _1534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5073__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_77_Left_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3703__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4820__A2 _2207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6599__CLK clknet_leaf_17_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5781__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5533__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3318__C _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5836__A1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3311__A2 _1055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput9 c0_o_instr_long_addr[4] net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3900_ _1384_ immu_0.page_table\[12\]\[5\] _1390_ _1565_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4880_ _1994_ _2241_ _2243_ net1004 _2256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6013__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3831_ _1368_ _1491_ _1497_ _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_39_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4575__A1 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3762_ _1372_ _1381_ _1430_ _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6550_ _0123_ clknet_leaf_6_core_clock immu_0.page_table\[6\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5772__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5501_ _2300_ _2629_ _2631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_82_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6481_ _0054_ clknet_leaf_33_core_clock dmmu0.page_table\[7\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3693_ _1350_ net311 _1360_ _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4327__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5432_ _2461_ _2582_ _2584_ net947 _2591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_83_core_clock_I clknet_4_10__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4878__A2 _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5363_ _2550_ _0222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7102_ net211 net517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4314_ _1915_ _0617_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5294_ _2510_ _0193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7033_ net288 net439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4245_ net198 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4176_ _1814_ _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3933__S0 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3127_ _0876_ _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_2_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input217_I dcache_mem_o_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3066__A1 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3058_ _0829_ net479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6741__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4263__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4802__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3161__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_2682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_2693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6817_ _0390_ clknet_leaf_67_core_clock dmmu1.page_table\[11\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6748_ _0321_ clknet_leaf_34_core_clock dmmu0.page_table\[6\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5763__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6679_ _0252_ clknet_leaf_37_core_clock dmmu0.page_table\[2\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5515__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_2486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_2497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5818__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output436_I net436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6271__CLK clknet_leaf_91_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3924__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output603_I net603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7140__I net389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3057__A1 net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_1309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6614__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_55_1858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4030_ immu_1.page_table\[12\]\[9\] immu_1.page_table\[13\]\[9\] immu_1.page_table\[14\]\[9\]
+ immu_1.page_table\[15\]\[9\] _1409_ _1410_ _1691_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5285__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Right_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4493__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7050__I net286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5037__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5981_ _1770_ _2906_ _2908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4932_ _2289_ _2292_ _1771_ _0049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3599__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5993__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4863_ _2247_ _0025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6602_ _0175_ clknet_leaf_8_core_clock immu_0.page_table\[2\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_14 net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3814_ _1434_ net705 _1476_ _1481_ _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA_25 net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4794_ _2171_ net76 _2205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_27_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6533_ _0106_ clknet_leaf_5_core_clock immu_0.page_table\[8\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3745_ net369 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_43_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6464_ _0037_ clknet_leaf_30_core_clock dmmu0.page_table\[8\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3676_ _1350_ net322 _1326_ _1351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5415_ _2580_ _0244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6294__CLK clknet_leaf_90_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6395_ _0777_ clknet_leaf_1_core_clock immu_0.page_table\[15\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4720__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input167_I c1_o_req_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5346_ _2455_ _2536_ _2538_ net782 _2542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_71_2350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5277_ _1776_ _2500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input334_I ic1_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4228_ _1857_ _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_78_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3287__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input28_I c0_o_mem_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4159_ net98 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_84_2733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_2154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_2176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4251__A3 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_2010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4539__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5736__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_inner_720 c1_i_core_int_sreg[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_68_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinterconnect_inner_731 c1_i_core_int_sreg[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_18_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5200__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_2548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6637__CLK clknet_leaf_11_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3762__A2 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output553_I net553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6161__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7135__I net65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6787__CLK clknet_leaf_44_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5267__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3278__A1 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3373__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3104__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5019__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4778__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 c0_o_instr_long_addr[7] net12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput23 c0_o_mem_addr[4] net23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput34 c0_o_mem_data[14] net34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput45 c0_o_mem_high_addr[0] net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3530_ _1264_ net551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4950__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4950__B2 dmmu0.page_table\[7\]\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput56 c0_o_mem_sel[1] net56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput67 c0_o_req_addr[2] net67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput78 c0_sr_bus_addr[11] net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput89 c0_sr_bus_addr[7] net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3461_ _0912_ _1195_ _1200_ _1201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7045__I net281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5200_ _2453_ _2447_ _2449_ immu_0.page_table\[3\]\[2\] _2454_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_27_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4702__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6180_ _3021_ _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3392_ dmmu1.page_table\[8\]\[8\] dmmu1.page_table\[9\]\[8\] dmmu1.page_table\[10\]\[8\]
+ dmmu1.page_table\[11\]\[8\] _0887_ _0909_ _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5131_ _2410_ _0130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5062_ _2371_ _0100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3269__A1 net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4013_ immu_0.page_table\[12\]\[8\] immu_0.page_table\[13\]\[8\] immu_0.page_table\[14\]\[8\]
+ immu_0.page_table\[15\]\[8\] _1487_ _1390_ _1675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3522__B _1259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5964_ _2898_ _0475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5430__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4915_ _1819_ _2261_ _2263_ net805 _2280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3441__A1 net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5895_ _2782_ _2856_ _2858_ net1030 _2860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5718__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4846_ _2236_ _0019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5194__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4777_ _2196_ _0799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input284_I ic0_mem_data[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6516_ _0089_ clknet_leaf_8_core_clock immu_0.page_table\[9\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3728_ _1385_ immu_0.page_table\[5\]\[0\] _1397_ _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_73_2401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6447_ _0020_ clknet_leaf_102_core_clock dmmu0.page_table\[10\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3659_ _1337_ net248 _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5497__A2 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6378_ _0760_ clknet_leaf_78_core_clock immu_1.page_table\[11\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5329_ net93 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_60_1868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5404__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4457__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_2238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4209__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3680__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5957__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_2059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3983__A2 _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_29_core_clock clknet_4_5__leaf_core_clock clknet_leaf_29_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_81_1058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4696__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4999__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3346__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3671__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6802__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Left_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_1094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3423__A1 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4700_ _2067_ _2139_ _2142_ net1085 _2149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5680_ _2063_ _2726_ _2728_ dmmu1.page_table\[13\]\[4\] _2733_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4631_ _2107_ _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_leaf_68_core_clock clknet_4_12__leaf_core_clock clknet_leaf_68_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5176__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5783__I _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_22_core_clock_I clknet_4_4__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4562_ _2066_ _0714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6301_ _0683_ clknet_leaf_88_core_clock immu_1.page_table\[1\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3513_ dmmu1.page_table\[0\]\[12\] dmmu1.page_table\[1\]\[12\] dmmu1.page_table\[2\]\[12\]
+ dmmu1.page_table\[3\]\[12\] _0886_ _0900_ _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_69_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4493_ _1858_ _2014_ _2016_ immu_1.page_table\[3\]\[5\] _2022_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5479__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6232_ _0614_ clknet_leaf_88_core_clock immu_1.page_table\[0\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_10__f_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_3444_ _1180_ _1183_ _1119_ _1184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3375_ _1114_ _1116_ _0879_ _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6163_ _2849_ _3000_ _3002_ net785 _3012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5114_ _2265_ _2398_ _2400_ immu_0.page_table\[6\]\[1\] _2402_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6094_ _2971_ _0532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4439__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5045_ _2275_ _2352_ _2354_ immu_0.page_table\[9\]\[6\] _2361_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3662__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Left_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6482__CLK clknet_leaf_32_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5939__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6996_ _0569_ clknet_leaf_97_core_clock dmmu1.long_off_reg\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_24_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3414__A1 net153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5947_ _2049_ _2872_ _2874_ net912 _2888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_24_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4611__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5878_ _2848_ _0439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input95_I c0_sr_bus_data_o[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_2079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4829_ _1797_ _2224_ _2226_ net1075 _2228_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3717__A2 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3427__B _1167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4678__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput202 c1_sr_bus_data_o[2] net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput213 dcache_mem_exception net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_60_1687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput224 dcache_mem_o_data[4] net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput235 dcache_wb_adr[13] net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput246 dcache_wb_adr[23] net246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput257 dcache_wb_o_dat[10] net257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput268 dcache_wb_o_dat[6] net268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output516_I net516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3328__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput279 ic0_mem_data[11] net279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5642__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3653__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6975__CLK clknet_leaf_105_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3500__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6205__CLK clknet_leaf_96_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4905__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6107__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4381__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6355__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_88_core_clock_I clknet_4_10__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4133__A2 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5330__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_2015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3160_ _0909_ _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_20_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3892__A1 net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold1 ic0_wb_cyc net735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_59_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3091_ net128 net23 _0842_ _0848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _0423_ clknet_leaf_39_core_clock dmmu0.page_table\[1\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5801_ _2805_ _0405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5397__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6781_ _0354_ clknet_leaf_47_core_clock dmmu1.page_table\[13\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_8_Right_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3993_ immu_1.page_table\[4\]\[8\] immu_1.page_table\[5\]\[8\] immu_1.page_table\[6\]\[8\]
+ immu_1.page_table\[7\]\[8\] _1404_ _1540_ _1655_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_85_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5732_ _2051_ _2760_ _2762_ net837 _2763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3947__A2 _1594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5149__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5663_ _2722_ _0350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4614_ _2097_ _0735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5594_ _2444_ _2681_ _2684_ net1078 _2685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4545_ _2054_ _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4476_ _2011_ _0683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6215_ _0597_ clknet_leaf_90_core_clock immu_1.page_table\[7\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4857__I _2243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5321__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4124__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3427_ _0912_ _1162_ _1167_ _0895_ _1168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XPHY_EDGE_ROW_39_Right_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input247_I dcache_wb_adr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5872__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6146_ _3003_ _0552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3358_ dmmu0.page_table\[8\]\[7\] dmmu0.page_table\[9\]\[7\] dmmu0.page_table\[10\]\[7\]
+ dmmu0.page_table\[11\]\[7\] _0950_ _0952_ _1101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_77_1436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6077_ _2784_ _2958_ _2960_ net784 _2963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3289_ dmmu0.page_table\[13\]\[4\] _1035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5085__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5624__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ _2350_ _0087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input10_I c0_o_instr_long_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3635__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6998__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_90_core_clock_I clknet_4_8__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5388__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6979_ _0552_ clknet_leaf_79_core_clock immu_1.page_table\[8\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_48_Right_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_1420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4060__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6378__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4899__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Right_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output633_I net633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7143__I net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_1981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_66_Right_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_1228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3485__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5551__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Right_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3788__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput506 net506 c1_i_req_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_2058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput517 net517 c1_rst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput528 net528 dcache_mem_addr[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4330_ _1923_ _0625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput539 net539 dcache_mem_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4106__A2 net327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ _1852_ _1876_ _1878_ net878 _1882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7053__I net290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6000_ _2918_ _0491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3212_ _0940_ _0883_ _0960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5854__A2 _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I c0_o_c_instr_long vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4192_ net188 _1827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__3865__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3143_ net124 _0892_ _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3960__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5067__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5606__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3074_ net219 _0831_ _0838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3617__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Right_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_2034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4814__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6902_ _0475_ clknet_leaf_57_core_clock dmmu1.page_table\[5\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6833_ _0406_ clknet_leaf_50_core_clock dmmu1.page_table\[9\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3957__S _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6031__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6764_ _0337_ clknet_leaf_34_core_clock dmmu0.page_table\[5\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3976_ _1637_ _1638_ _1366_ _1639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5715_ _2752_ _0372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4593__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5790__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6695_ _0268_ clknet_leaf_35_core_clock dmmu0.page_table\[4\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_1096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input197_I c1_sr_bus_data_o[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5646_ net94 _2698_ _2700_ net1056 _2713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_85_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3228__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3779__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5577_ _2069_ _2664_ _2666_ dmmu1.page_table\[15\]\[7\] _2674_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6670__CLK clknet_leaf_103_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold220 immu_1.page_table\[8\]\[1\] net954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input364_I ic1_wb_adr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold231 immu_0.page_table\[15\]\[7\] net965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4528_ _2043_ _0703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_83_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold242 immu_0.page_table\[11\]\[4\] net976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold253 immu_1.page_table\[15\]\[6\] net987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input58_I c0_o_req_active vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold264 immu_0.page_table\[2\]\[10\] net998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold275 dmmu0.page_table\[1\]\[3\] net1009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold286 immu_0.page_table\[13\]\[8\] net1020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4459_ _1845_ _1999_ _2001_ immu_1.page_table\[1\]\[1\] _2003_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xhold297 immu_1.page_table\[8\]\[7\] net1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7178_ net397 net650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6129_ net213 net212 _2991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5412__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3608__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3703__S1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5211__I _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4033__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5230__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output583_I net583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5781__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3219__S0 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5533__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5297__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5836__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5049__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6543__CLK clknet_leaf_23_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6013__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3830_ _1378_ _1381_ _1496_ _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4024__A1 net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3458__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5772__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3761_ _1368_ _1429_ _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4575__A2 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7048__I net284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6693__CLK clknet_leaf_91_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5500_ _2629_ _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_54_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6480_ _0053_ clknet_leaf_34_core_clock dmmu0.page_table\[7\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3692_ _1348_ net365 _1363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5431_ _2590_ _0250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4327__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5362_ _1994_ _2535_ _2537_ dmmu0.page_table\[15\]\[11\] _2550_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_65_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7101_ net330 net516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4313_ _1824_ _1911_ _1914_ immu_1.page_table\[2\]\[0\] _1915_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5293_ _1811_ _2502_ _2504_ immu_0.page_table\[0\]\[6\] _2510_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7032_ net277 net428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4244_ _1869_ _0593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3838__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4175_ net102 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3933__S1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3126_ _0875_ _0876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3260__B _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3057_ net226 _0822_ _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4263__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3066__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input112_I c1_o_instr_long_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_2683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6816_ _0389_ clknet_leaf_69_core_clock dmmu1.page_table\[11\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4015__A1 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5212__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6747_ _0320_ clknet_leaf_35_core_clock dmmu0.page_table\[6\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5763__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3959_ _1434_ _1621_ _1622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6678_ _0251_ clknet_leaf_40_core_clock dmmu0.page_table\[2\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_4_8__f_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5629_ _2704_ _0334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5515__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_2487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_2498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5818__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3829__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output429_I net429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3924__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6566__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3057__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_2057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5876__I net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5203__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5754__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3860__S0 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_27_core_clock_I clknet_4_5__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_2006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__CLK clknet_leaf_64_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4493__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5690__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3540__I0 net147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5980_ _2906_ _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_56_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5442__B1 _2583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4931_ _1776_ _2290_ _2291_ _1823_ _2292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5993__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4862_ _1800_ _2242_ _2244_ dmmu0.page_table\[9\]\[2\] _2247_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6601_ _0174_ clknet_leaf_19_core_clock immu_0.page_table\[2\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3813_ _1433_ _1477_ _1480_ _1415_ _1481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA_15 net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _2204_ _0807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_26 net404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6532_ _0105_ clknet_leaf_6_core_clock immu_0.page_table\[8\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3744_ immu_1.page_table\[12\]\[0\] immu_1.page_table\[13\]\[0\] immu_1.page_table\[14\]\[0\]
+ immu_1.page_table\[15\]\[0\] _1409_ _1410_ _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_12_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _0036_ clknet_leaf_30_core_clock dmmu0.page_table\[8\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3675_ _0813_ _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6439__CLK clknet_leaf_17_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5414_ immu_0.high_addr_off\[7\] _1815_ _2572_ _2580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6394_ _0776_ clknet_leaf_1_core_clock immu_0.page_table\[15\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5345_ _2541_ _0213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4720__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_2340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_2362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5276_ _2499_ _0186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6589__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4227_ net205 _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_78_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3531__I0 net143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input327_I ic0_wb_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4158_ _1801_ _0575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_1946 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_2734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3109_ net19 _0858_ _0859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_84_2745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ net116 immu_1.high_addr_off\[6\] _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_1269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_2177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_2033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinterconnect_inner_710 c0_i_core_int_sreg[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_inner_721 c1_i_core_int_sreg[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_80_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_inner_732 c1_i_core_int_sreg[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_18_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_2549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_19_core_clock clknet_4_4__leaf_core_clock clknet_leaf_19_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6161__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7151__I net391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__A1 net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5672__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5424__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4778__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5975__A1 net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_58_core_clock clknet_4_14__leaf_core_clock clknet_leaf_58_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_64_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 c0_o_mem_addr[0] net13 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3833__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput24 c0_o_mem_addr[5] net24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput35 c0_o_mem_data[15] net35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput46 c0_o_mem_high_addr[1] net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_29_1525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4950__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput57 c0_o_mem_we net57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput68 c0_o_req_addr[3] net68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput79 c0_sr_bus_addr[12] net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3460_ net123 _1197_ _1199_ _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_46_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6731__CLK clknet_leaf_100_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4702__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3790__S _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3391_ _0896_ _1132_ _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5130_ _2330_ _2398_ _2400_ net970 _2410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_1146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4685__I _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5061_ _2265_ _2367_ _2369_ immu_0.page_table\[8\]\[1\] _2371_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6881__CLK clknet_leaf_67_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4012_ _1367_ _1673_ _1674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_97_core_clock clknet_4_9__leaf_core_clock clknet_leaf_97_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_7_1928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5963_ _2790_ _2890_ _2892_ dmmu1.page_table\[5\]\[5\] _2898_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4914_ _2279_ _0044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5894_ _2859_ _0444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_95_core_clock_I clknet_4_8__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_2030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4845_ _1819_ _2224_ _2226_ net758 _2236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5718__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6261__CLK clknet_leaf_85_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4776_ _1800_ _2191_ _2193_ immu_0.page_table\[12\]\[2\] _2196_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5194__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3824__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6515_ _0088_ clknet_leaf_3_core_clock immu_0.page_table\[9\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3727_ _1396_ immu_0.page_table\[4\]\[0\] _1397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3764__I _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_2413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input277_I ic0_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6143__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6446_ _0019_ clknet_leaf_15_core_clock dmmu0.page_table\[10\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3658_ inner_wb_arbiter.o_sel_sig _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_30_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6377_ _0759_ clknet_leaf_74_core_clock immu_1.page_table\[11\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3589_ net216 _1219_ _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5328_ _2530_ _0207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input40_I c0_o_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5259_ _1799_ _2486_ _2488_ immu_0.page_table\[1\]\[2\] _2491_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4457__A1 _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_2217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4209__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3680__A2 net323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5957__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6604__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output496_I net496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3196__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7146__I net401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_2101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_1910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4696__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5893__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_33_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4448__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4999__A2 _2316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3671__A2 net251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6284__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3785__S _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4059__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4630_ _1838_ _1892_ _2028_ _2107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_56_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5176__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_2012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4561_ _2065_ _2053_ _2055_ net779 _2066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7056__I net293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6300_ _0682_ clknet_leaf_88_core_clock immu_1.page_table\[1\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_1847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3512_ net157 dmmu1.long_off_reg\[7\] _1249_ _1250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_40_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6125__A1 net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4492_ _2021_ _0689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6231_ _0613_ clknet_leaf_85_core_clock immu_1.page_table\[0\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3443_ _1142_ _1181_ _1182_ _1183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_46_1691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6162_ _3011_ _0560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3374_ _0940_ _1115_ _1116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5113_ _2401_ _0121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_85_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6093_ _2851_ _2957_ _2959_ dmmu1.page_table\[1\]\[10\] _2971_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5304__I _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4439__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5636__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5044_ _2360_ _0093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3252__C _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3111__A1 net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6627__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_2049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3662__A2 net319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5939__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6995_ _0568_ clknet_leaf_97_core_clock dmmu1.long_off_reg\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6061__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ _2887_ _0468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4611__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6777__CLK clknet_leaf_103_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5877_ _2847_ _2836_ _2838_ dmmu1.page_table\[8\]\[8\] _2848_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_79_2600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input394_I inner_wb_i_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4828_ _2227_ _0010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4375__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input88_I c0_sr_bus_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4759_ _1815_ _2175_ _2177_ net746 _2185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3427__C _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6429_ _0002_ clknet_leaf_110_core_clock immu_0.page_table\[13\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4678__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_8_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3350__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput203 c1_sr_bus_data_o[3] net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_1065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput214 dcache_mem_o_data[0] net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput225 dcache_mem_o_data[5] net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5214__I _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput236 dcache_wb_adr[14] net236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput247 dcache_wb_adr[2] net247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput258 dcache_wb_o_dat[11] net258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput269 dcache_wb_o_dat[7] net269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output509_I net509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3653__A2 net317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_9_core_clock clknet_4_1__leaf_core_clock clknet_leaf_9_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3169__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4905__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6107__A1 _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5866__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5330__A2 _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_105_core_clock clknet_4_2__leaf_core_clock clknet_leaf_105_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_24_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold2 immu_1.page_table\[0\]\[0\] net736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3090_ _0847_ net535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4841__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6043__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5800_ _2776_ _2802_ _2804_ net1023 _2805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_18_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6780_ _0353_ clknet_leaf_47_core_clock dmmu1.page_table\[13\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3992_ _1651_ _1652_ _1653_ _1654_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5397__A2 net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5731_ _2761_ _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_15_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5662_ dmmu0.long_off_reg\[5\] _1809_ _2716_ _2722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5149__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4357__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4613_ _2063_ _2090_ _2092_ immu_1.page_table\[13\]\[4\] _2097_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5593_ _2683_ _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_13_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4544_ _1912_ _2052_ _2054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3247__C _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4475_ net209 _1999_ _2001_ immu_1.page_table\[1\]\[9\] _2011_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_1_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_2042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6214_ _0596_ clknet_leaf_87_core_clock immu_1.page_table\[7\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3426_ _1164_ _1166_ net123 _1167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__5321__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6145_ _1823_ _3000_ _3002_ immu_1.page_table\[8\]\[0\] _3003_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3357_ _0940_ _1099_ _1100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input142_I c1_o_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6076_ _2962_ _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3288_ _0882_ _1032_ _1033_ _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_1448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5085__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _2332_ _2336_ _2338_ net1011 _2350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3635__A2 net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4094__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_2111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5388__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6978_ _0551_ clknet_leaf_105_core_clock mem_dcache_arb.transfer_active vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3238__I2 dmmu1.page_table\[14\]\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3399__A1 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_1481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5929_ _2786_ _2873_ _2875_ net745 _2879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4899__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3571__A1 net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output459_I net459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5848__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5879__I net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6942__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3901__B _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6025__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4587__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3485__S1 _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6179__I1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6322__CLK clknet_leaf_70_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4339__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5551__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_2037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput507 net507 c1_i_req_data[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput518 net518 dcache_mem_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput529 net529 dcache_mem_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6472__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4260_ _1881_ _0597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3211_ _0956_ _0957_ _0958_ _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4191_ net190 _1825_ _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_24_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3142_ _0890_ _0891_ _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5067__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3073_ _0837_ net471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4814__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3617__A2 net265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3173__S0 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6901_ _0474_ clknet_leaf_53_core_clock dmmu1.page_table\[5\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_34_core_clock_I clknet_4_7__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _0405_ clknet_leaf_50_core_clock dmmu1.page_table\[9\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6763_ _0336_ clknet_leaf_37_core_clock dmmu0.page_table\[5\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3975_ immu_0.page_table\[4\]\[7\] immu_0.page_table\[5\]\[7\] immu_0.page_table\[6\]\[7\]
+ immu_0.page_table\[7\]\[7\] _1396_ _1371_ _1638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_11_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5714_ _2067_ _2743_ _2745_ net926 _2752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6694_ _0267_ clknet_leaf_34_core_clock dmmu0.page_table\[4\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5645_ _2712_ _0342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3228__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6815__CLK clknet_leaf_44_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_2115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5576_ _2673_ _0312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold210 dmmu1.page_table\[4\]\[0\] net944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4527_ _1864_ _2033_ _2035_ dmmu1.page_table\[14\]\[7\] _2043_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold221 dmmu1.page_table\[3\]\[9\] net955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3772__I net366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold232 immu_0.page_table\[4\]\[6\] net966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold243 immu_0.page_table\[7\]\[10\] net977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold254 dmmu1.page_table\[4\]\[2\] net988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input357_I ic1_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold265 dmmu1.page_table\[3\]\[8\] net999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold276 immu_1.page_table\[2\]\[5\] net1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4458_ _2002_ _0674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold287 dmmu1.page_table\[2\]\[10\] net1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6965__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3305__A1 net150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold298 immu_1.page_table\[11\]\[6\] net1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_22_1734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3409_ dmmu0.page_table\[0\]\[9\] dmmu0.page_table\[1\]\[9\] dmmu0.page_table\[2\]\[9\]
+ dmmu0.page_table\[3\]\[9\] _0863_ _0866_ _1150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7177_ net396 net649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4389_ _1912_ _1956_ _1958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6128_ _2990_ _0547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6059_ _2847_ _2941_ _2943_ dmmu1.page_table\[2\]\[8\] _2952_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3608__A2 net274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6345__CLK clknet_leaf_63_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4569__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5230__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5781__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6495__CLK clknet_leaf_32_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3219__S1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5533__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7154__I net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_2092 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5297__A1 net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5049__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_2052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5221__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3458__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3083__I0 net118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3760_ immu_0.page_table\[2\]\[1\] immu_0.page_table\[3\]\[1\] immu_0.page_table\[10\]\[1\]
+ immu_0.page_table\[11\]\[1\] _1424_ _1377_ _1429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_27_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5772__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4575__A3 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3783__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3691_ _1359_ _1361_ _1362_ net661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3793__S _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5430_ _2459_ _2582_ _2584_ net992 _2590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_49_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6988__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4732__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5361_ _2549_ _0221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7100_ net355 net508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4312_ _1913_ _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5292_ _2509_ _0192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_1789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7031_ net406 net409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6218__CLK clknet_leaf_90_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4243_ _1868_ _1841_ _1843_ immu_1.page_table\[9\]\[9\] _1869_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4174_ _1813_ _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3125_ net17 _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6368__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3056_ _0828_ net478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4263__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input105_I c0_sr_bus_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_2673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_2684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ _0388_ clknet_leaf_44_core_clock dmmu1.page_table\[11\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5212__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6746_ _0319_ clknet_leaf_32_core_clock dmmu0.page_table\[6\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5763__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3958_ immu_1.page_table\[12\]\[7\] immu_1.page_table\[13\]\[7\] immu_1.page_table\[14\]\[7\]
+ immu_1.page_table\[15\]\[7\] _1441_ _1442_ _1621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_73_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3889_ net6 immu_0.high_addr_off\[1\] _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6677_ _0250_ clknet_leaf_38_core_clock dmmu0.page_table\[2\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5628_ _1799_ _2699_ _2701_ net786 _2704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5515__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input70_I c0_o_req_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_2488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5559_ _1874_ _2028_ _2031_ _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_76_2499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5451__A1 _1834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3462__B1 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5203__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_48_core_clock clknet_4_13__leaf_core_clock clknet_leaf_48_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7149__I net404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_2_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4962__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3860__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3517__A1 _0905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_2018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_1974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6510__CLK clknet_leaf_6_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4493__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5690__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3540__I1 net42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_87_core_clock clknet_4_10__leaf_core_clock clknet_leaf_87_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_63_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5442__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4971__I _2316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4930_ _1829_ _1837_ _2286_ _2291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__6660__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5993__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4861_ _2246_ _0024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6600_ _0173_ clknet_leaf_22_core_clock immu_0.page_table\[2\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3812_ _1433_ _1478_ _1479_ _1480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_7_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4792_ _1821_ _2190_ _2192_ immu_0.page_table\[12\]\[10\] _2204_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_16 net396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_27 net404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3300__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3743_ immu_1.page_table\[4\]\[0\] immu_1.page_table\[5\]\[0\] immu_1.page_table\[6\]\[0\]
+ immu_1.page_table\[7\]\[0\] _1409_ _1410_ _1413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6531_ _0104_ clknet_leaf_4_core_clock immu_0.page_table\[8\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6462_ _0035_ clknet_leaf_103_core_clock dmmu0.page_table\[9\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3674_ _1348_ net376 _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3508__A1 _1119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5413_ _2579_ _0243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6393_ _0775_ clknet_leaf_109_core_clock immu_0.page_table\[15\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5344_ _2453_ _2536_ _2538_ net885 _2541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_71_2341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_2352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5275_ net93 _2485_ _2487_ immu_0.page_table\[1\]\[10\] _2499_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_80_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4226_ _1856_ _0588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5130__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3531__I1 net38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4157_ _1800_ _1792_ _1794_ net1028 _1801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input222_I dcache_mem_o_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3119__S0 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3108_ _0856_ _0857_ _0858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_84_2724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_2735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4088_ _1350_ _1579_ _1746_ _1747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_84_2746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3039_ mem_dcache_arb.select _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_65_2156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_65_2178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5197__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5736__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_inner_711 c0_i_core_int_sreg[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_18_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinterconnect_inner_722 c1_i_core_int_sreg[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_19_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_inner_733 c1_i_core_int_sreg[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4944__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6729_ _0302_ clknet_leaf_14_core_clock dmmu0.page_table\[3\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_22_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_22_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6161__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6533__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output441_I net441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput690 net690 inner_wb_o_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3358__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3181__B _0929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5672__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_6_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6683__CLK clknet_leaf_101_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5424__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5975__A2 _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_1653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_1664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4935__B1 _2291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 c0_o_mem_addr[10] net14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3833__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput25 c0_o_mem_addr[6] net25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput36 c0_o_mem_data[1] net36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput47 c0_o_mem_high_addr[2] net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput58 c0_o_req_active net58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput69 c0_o_req_addr[4] net69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3390_ dmmu1.page_table\[12\]\[8\] dmmu1.page_table\[13\]\[8\] dmmu1.page_table\[14\]\[8\]
+ dmmu1.page_table\[15\]\[8\] _0887_ _0909_ _1132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_0_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3910__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_15__f_core_clock clknet_3_7_0_core_clock clknet_4_15__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_23_1158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5060_ _2370_ _0099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5112__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4011_ immu_0.page_table\[8\]\[8\] immu_0.page_table\[9\]\[8\] immu_0.page_table\[10\]\[8\]
+ immu_0.page_table\[11\]\[8\] _1487_ _1390_ _1673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_74_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5962_ _2897_ _0474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4913_ _1817_ _2261_ _2263_ dmmu0.page_table\[8\]\[8\] _2279_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5893_ _2776_ _2856_ _2858_ net891 _2859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_60_2020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_2031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5718__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4844_ _2235_ _0018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_16_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3729__B2 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4775_ _2195_ _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3824__S1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6514_ _0087_ clknet_leaf_2_core_clock immu_0.page_table\[10\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3726_ _1369_ _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_28_1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6556__CLK clknet_leaf_23_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_73_2403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6445_ _0018_ clknet_leaf_26_core_clock dmmu0.page_table\[10\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_2414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3657_ _0814_ net318 _1326_ _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input172_I c1_o_req_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3588_ _1294_ net412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6376_ _0758_ clknet_leaf_75_core_clock immu_1.page_table\[11\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5327_ _2529_ _2516_ _2518_ dmmu0.page_table\[12\]\[9\] _2530_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5103__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5258_ _2490_ _0177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input33_I c0_o_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4457__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4209_ _1824_ _1841_ _1843_ immu_1.page_table\[9\]\[0\] _1844_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5189_ _1780_ _1971_ _2445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_67_2218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3760__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4209__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5957__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3221__S _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5500__I _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_2006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4116__I _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4917__B1 _2262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output489_I net489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_1900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5342__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5893__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4696__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7162__I net176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4448__A2 _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6429__CLK clknet_leaf_110_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3959__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_39_core_clock_I clknet_4_6__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4059__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6579__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4908__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4560_ _1857_ _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_25_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5581__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3511_ _1216_ _1247_ _1248_ _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4491_ _1855_ _2014_ _2016_ net1053 _2021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6125__A2 _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3442_ net49 dmmu0.long_off_reg\[4\] _1182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6230_ _0612_ clknet_leaf_82_core_clock immu_1.page_table\[0\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3373_ dmmu0.page_table\[4\]\[8\] dmmu0.page_table\[5\]\[8\] dmmu0.page_table\[6\]\[8\]
+ dmmu0.page_table\[7\]\[8\] _0864_ _0941_ _1115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6161_ _2847_ _3000_ _3002_ net908 _3011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7072__I net356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5112_ _2258_ _2398_ _2400_ immu_0.page_table\[6\]\[0\] _2401_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6092_ _2970_ _0531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5636__A1 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4439__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5043_ _2273_ _2352_ _2354_ immu_0.page_table\[9\]\[5\] _2360_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3105__I _0855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3111__A2 net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3742__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6994_ _0567_ clknet_leaf_97_core_clock dmmu1.long_off_reg\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5939__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6061__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5945_ _2047_ _2872_ _2874_ net879 _2887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_2004 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4611__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3976__S _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5876_ net208 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_5_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_2601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4827_ _1777_ _2224_ _2226_ net888 _2227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input387_I inner_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4375__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4758_ _2184_ _0792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_1412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3709_ _1375_ _1376_ _1378_ _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_31_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4689_ _2143_ _0764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4127__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5324__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6428_ _0001_ clknet_leaf_110_core_clock immu_0.page_table\[13\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_41_core_clock_I clknet_4_6__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4678__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6359_ _0741_ clknet_leaf_71_core_clock immu_1.page_table\[13\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3216__S _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput204 c1_sr_bus_data_o[4] net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3350__A2 _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput215 dcache_mem_o_data[10] net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput226 dcache_mem_o_data[6] net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_1088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput237 dcache_wb_adr[15] net237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput248 dcache_wb_adr[3] net248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput259 dcache_wb_o_dat[12] net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_58_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6721__CLK clknet_leaf_41_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7157__I net171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5402__I1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6871__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5563__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6107__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5315__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5866__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_1128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5618__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6251__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold3 immu_0.page_table\[0\]\[0\] net737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_55_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4841__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_2050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6043__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3991_ _1651_ _1652_ net107 _1653_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5730_ _2682_ _2759_ _2761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_50_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5661_ _2721_ _0349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7067__I net407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4357__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4612_ _2096_ _0734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_83_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5592_ _2682_ _2680_ _2683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_26_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ _2052_ _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4109__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4474_ _2010_ _0682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6213_ _0595_ clknet_leaf_84_core_clock immu_1.page_table\[7\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3425_ _0906_ _1165_ _1166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_2076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3356_ dmmu0.page_table\[12\]\[7\] dmmu0.page_table\[13\]\[7\] dmmu0.page_table\[14\]\[7\]
+ dmmu0.page_table\[15\]\[7\] _0882_ _0948_ _1099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6144_ _3001_ _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_42_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3287_ _0882_ dmmu0.page_table\[14\]\[4\] _0941_ _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6075_ _2782_ _2958_ _2960_ net1006 _2962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5085__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input135_I c1_o_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5026_ _2349_ _0086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6744__CLK clknet_leaf_69_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4293__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3486__I3 dmmu0.page_table\[3\]\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input302_I ic0_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4045__B1 _1705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6977_ _0550_ clknet_leaf_105_core_clock mem_dcache_arb.req0_pending vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5928_ _2878_ _0459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6894__CLK clknet_leaf_67_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5859_ _2837_ _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_64_958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5545__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4899__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3571__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5848__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6274__CLK clknet_leaf_89_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5225__I _2469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output521_I net521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3706__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4823__A2 _2222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6025__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4587__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5784__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4339__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_3__f_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6617__CLK clknet_leaf_24_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_2049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput508 net508 c1_i_req_data[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_50_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput519 net519 dcache_mem_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3210_ net18 _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__4511__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4190_ net189 _1825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__6767__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3141_ net151 net150 net153 net152 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_EDGE_ROW_19_Left_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5067__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3072_ net218 _0831_ _0837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_2014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4814__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6900_ _0473_ clknet_leaf_55_core_clock dmmu1.page_table\[5\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3173__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_2058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6831_ _0404_ clknet_leaf_68_core_clock dmmu1.page_table\[10\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5775__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6762_ _0335_ clknet_leaf_48_core_clock dmmu0.page_table\[5\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_1898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3974_ immu_0.page_table\[0\]\[7\] immu_0.page_table\[1\]\[7\] immu_0.page_table\[2\]\[7\]
+ immu_0.page_table\[3\]\[7\] _1396_ _1371_ _1637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_50_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5713_ _2751_ _0371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6693_ _0266_ clknet_leaf_91_core_clock immu_1.high_addr_off\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_28_Left_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_1076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_2110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3258__C _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5527__B1 _2631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5644_ _2531_ _2698_ _2700_ net1041 _2712_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6297__CLK clknet_leaf_82_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5575_ _2067_ _2664_ _2666_ dmmu1.page_table\[15\]\[6\] _2673_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_83_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold200 immu_1.page_table\[2\]\[2\] net934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_25_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold211 immu_1.page_table\[6\]\[6\] net945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4526_ _2042_ _0702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold222 immu_0.page_table\[8\]\[8\] net956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_14_899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold233 immu_1.page_table\[6\]\[5\] net967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold244 immu_1.page_table\[14\]\[6\] net978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold255 dmmu1.page_table\[7\]\[2\] net989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4457_ _1823_ _1999_ _2001_ immu_1.page_table\[1\]\[0\] _2002_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xhold266 dmmu0.page_table\[2\]\[0\] net1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold277 immu_0.page_table\[10\]\[10\] net1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input252_I dcache_wb_adr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold288 immu_0.page_table\[5\]\[7\] net1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold299 immu_1.page_table\[4\]\[4\] net1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_22_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3936__S0 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3408_ _0875_ _1148_ _1149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7176_ net389 net642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4388_ _1956_ _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_37_Left_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4884__I _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6127_ net200 _2974_ _2976_ dmmu1.page_table\[0\]\[12\] _2990_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3339_ _1069_ _1080_ _1081_ _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_77_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _2951_ _0516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5009_ _2265_ _2337_ _2339_ immu_0.page_table\[10\]\[1\] _2341_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6007__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4018__B1 _1669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4569__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_38_core_clock clknet_4_6__leaf_core_clock clknet_leaf_38_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5766__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Left_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5230__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3241__A1 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5297__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Left_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_53_1799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5049__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_77_core_clock clknet_4_11__leaf_core_clock clknet_leaf_77_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4257__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_64_Left_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5221__A2 _2446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3359__B _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5509__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3690_ _1337_ net232 _1362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4732__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5360_ _2531_ _2535_ _2537_ net937 _2549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4311_ _1912_ _1910_ _1913_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5291_ _1808_ _2502_ _2504_ immu_0.page_table\[0\]\[5\] _2509_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7030_ net386 net408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4242_ net209 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3299__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4173_ _1812_ _1792_ _1794_ immu_0.page_table\[11\]\[6\] _1813_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7080__I net333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3124_ dmmu0.page_table\[8\]\[0\] dmmu0.page_table\[9\]\[0\] dmmu0.page_table\[10\]\[0\]
+ dmmu0.page_table\[11\]\[0\] _0872_ _0868_ _0874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_74_1419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3055_ net225 _0822_ _0828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3113__I net15 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_2674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6814_ _0387_ clknet_leaf_45_core_clock dmmu1.page_table\[11\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5748__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5212__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3223__A1 _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6745_ _0318_ clknet_leaf_69_core_clock dmmu1.page_table\[15\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3957_ _1618_ _1619_ _1416_ _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6676_ _0249_ clknet_leaf_38_core_clock dmmu0.page_table\[2\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3888_ net5 immu_0.high_addr_off\[0\] _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_34_939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5627_ _2703_ _0333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6932__CLK clknet_leaf_62_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5558_ _2662_ _0305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_76_2489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input63_I c0_o_req_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4509_ _1909_ _2028_ _2031_ _2032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5489_ _2527_ _2613_ _2615_ dmmu0.page_table\[4\]\[8\] _2624_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4487__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7159_ net173 net629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6312__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5987__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3462__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3462__B2 _1201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6462__CLK clknet_leaf_103_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5203__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3907__B _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7165__I net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4714__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5911__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5690__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6805__CLK clknet_leaf_69_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5442__A2 _2581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4650__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4860_ _1797_ _2242_ _2244_ dmmu0.page_table\[9\]\[1\] _2246_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3811_ _1474_ immu_1.page_table\[15\]\[2\] _1479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6955__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4791_ _2203_ _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_83_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_17 net396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_28 _1262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6530_ _0103_ clknet_leaf_3_core_clock immu_0.page_table\[8\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3742_ immu_1.page_table\[8\]\[0\] immu_1.page_table\[9\]\[0\] immu_1.page_table\[10\]\[0\]
+ immu_1.page_table\[11\]\[0\] _1409_ _1410_ _1412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_43_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3300__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6155__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6461_ _0034_ clknet_leaf_13_core_clock dmmu0.page_table\[9\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3673_ _1301_ _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7075__I net359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5412_ immu_0.high_addr_off\[6\] _1812_ _2572_ _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_1109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6392_ _0774_ clknet_leaf_98_core_clock immu_1.page_table\[10\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5343_ _2540_ _0212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_2342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_71_2353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_46_core_clock_I clknet_4_13__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6335__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5274_ _2498_ _0185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4469__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4225_ _1855_ _1841_ _1843_ immu_1.page_table\[9\]\[4\] _1856_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5130__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5323__I net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4156_ _1799_ _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_39_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3692__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6485__CLK clknet_leaf_32_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3119__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3107_ net46 net45 net48 net47 _0857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_TAPCELL_ROW_84_2725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5969__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4087_ net12 immu_0.high_addr_off\[7\] _1745_ _1746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA_input215_I dcache_mem_o_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3038_ _0812_ _0814_ _0816_ net603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_17_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_2157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_2168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_2179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_2057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5197__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4989_ _2327_ _0071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinterconnect_inner_712 c0_i_core_int_sreg[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_inner_723 c1_i_core_int_sreg[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4944__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6728_ _0301_ clknet_leaf_44_core_clock dmmu0.page_table\[3\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinterconnect_inner_734 c1_i_irq vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_22_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_2057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6659_ _0232_ clknet_leaf_26_core_clock dmmu0.page_table\[11\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_4__f_core_clock clknet_3_2_0_core_clock clknet_4_4__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_30_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput680 net680 inner_wb_adr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput691 net691 inner_wb_o_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_79_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output434_I net434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_2085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3358__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6828__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3181__C _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5672__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3683__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4880__B1 _2243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5424__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6978__CLK clknet_leaf_105_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3435__A1 _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3986__A2 _1647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6208__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4935__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4935__B2 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput15 c0_o_mem_addr[11] net15 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput26 c0_o_mem_addr[7] net26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput37 c0_o_mem_data[2] net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput48 c0_o_mem_high_addr[3] net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput59 c0_o_req_addr[0] net59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_1798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6358__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5360__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3910__A2 _1560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5112__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4010_ _1670_ _1671_ _1367_ _1672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3674__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6175__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5961_ _2788_ _2890_ _2892_ dmmu1.page_table\[5\]\[4\] _2897_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4912_ _2278_ _0043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_1282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5892_ _2857_ _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_59_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_2010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_2019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_2021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4843_ _1817_ _2224_ _2226_ dmmu0.page_table\[10\]\[8\] _2235_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4774_ _1797_ _2191_ _2193_ immu_0.page_table\[12\]\[1\] _2195_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6513_ _0086_ clknet_leaf_5_core_clock immu_0.page_table\[10\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3725_ _1370_ immu_0.page_table\[6\]\[0\] _1391_ _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_2540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6444_ _0017_ clknet_leaf_25_core_clock dmmu0.page_table\[10\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_2404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3656_ _1302_ net372 _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_73_2415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6375_ _0757_ clknet_leaf_80_core_clock immu_1.page_table\[11\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3587_ net215 _1219_ _1294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input165_I c1_o_req_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5326_ net104 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_3_2_0_core_clock clknet_0_core_clock clknet_3_2_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_80_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5103__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5257_ _1796_ _2486_ _2488_ immu_0.page_table\[1\]\[1\] _2490_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_input332_I ic1_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4208_ _1842_ _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_3_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3665__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5188_ _1776_ _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_input26_I c0_o_mem_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4862__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4892__I _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_2219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4139_ net90 _1782_ _1784_ _1785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_19_1718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3760__S1 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3417__A1 net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4090__A1 net117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4917__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6500__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6119__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4132__I net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5342__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5893__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3656__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3408__A1 _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4605__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4081__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4908__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5581__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_2058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3510_ net156 dmmu1.long_off_reg\[6\] _1248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4490_ _2020_ _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3441_ net49 dmmu0.long_off_reg\[4\] _1181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6160_ _3010_ _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_1584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3372_ _0938_ _1113_ _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5111_ _2399_ _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6091_ _2849_ _2958_ _2960_ net778 _2970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5097__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5636__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5042_ _2359_ _0092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_1281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3742__S1 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6993_ _0566_ clknet_leaf_94_core_clock dmmu1.long_off_reg\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6061__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3121__I _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5944_ _2886_ _0467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4072__A1 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6523__CLK clknet_leaf_6_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5875_ _2846_ _0438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_2049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_2602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4826_ _2225_ _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_63_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5021__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4375__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4757_ _1812_ _2175_ _2177_ net762 _2184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6673__CLK clknet_leaf_41_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input282_I ic0_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3708_ _1377_ _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_71_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4688_ _2051_ _2139_ _2142_ net880 _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5324__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6427_ _0000_ clknet_leaf_108_core_clock immu_0.page_table\[13\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4127__A2 _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4887__I _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3639_ _0812_ net261 _1323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3335__B1 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6358_ _0740_ clknet_leaf_78_core_clock immu_1.page_table\[13\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3886__A1 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_8_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5309_ _2451_ _2516_ _2518_ net853 _2520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput205 c1_sr_bus_data_o[5] net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6289_ _0671_ clknet_leaf_100_core_clock dmmu0.page_table\[0\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput216 dcache_mem_o_data[11] net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput227 dcache_mem_o_data[7] net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput238 dcache_wb_adr[16] net238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput249 dcache_wb_adr[4] net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4835__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4063__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output599_I net599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5563__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5315__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4797__I _2207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7173__I net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5866__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3877__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_2007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5618__A2 _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3629__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold4 icore_sregs.c1_disable net738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_55_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6043__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_18_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3990_ net114 immu_1.high_addr_off\[4\] _1652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_18_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ dmmu0.long_off_reg\[4\] _1806_ _2716_ _2721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_84_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4611_ _2061_ _2090_ _2092_ immu_1.page_table\[13\]\[3\] _2096_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4357__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5591_ _1769_ _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_48_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4542_ _1838_ _1874_ _2028_ _2052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_40_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4109__A2 net255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4473_ net208 _1999_ _2001_ immu_1.page_table\[1\]\[8\] _2010_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7083__I net336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6212_ _0594_ clknet_leaf_97_core_clock immu_1.page_table\[9\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3424_ dmmu1.page_table\[0\]\[9\] dmmu1.page_table\[1\]\[9\] dmmu1.page_table\[2\]\[9\]
+ dmmu1.page_table\[3\]\[9\] _0886_ _0900_ _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_61_1944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3868__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3868__B2 net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6143_ _1980_ _2999_ _3001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3355_ _0938_ _1097_ _0879_ _1098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3116__I net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6074_ _2961_ _0522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3286_ dmmu0.page_table\[15\]\[4\] _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_13_Left_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5025_ _2330_ _2337_ _2339_ net1094 _2349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4293__A1 _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input128_I c1_o_mem_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_28_core_clock clknet_4_5__leaf_core_clock clknet_leaf_28_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4045__A1 net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4045__B2 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6976_ _0549_ clknet_leaf_105_core_clock mem_dcache_arb.req1_pending vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5242__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5927_ _2784_ _2873_ _2875_ dmmu1.page_table\[6\]\[2\] _2878_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_49_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5858_ _2682_ _2835_ _2837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input93_I c0_sr_bus_data_o[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4809_ _2215_ _0003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5545__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_17_Right_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_1167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5789_ _2797_ _0401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5848__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3859__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6569__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Right_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_67_core_clock clknet_4_12__leaf_core_clock clknet_leaf_67_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4808__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output514_I net514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3706__S1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5481__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6025__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4036__A1 net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4587__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5784__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7168__I net167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4339__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_2077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3645__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput509 net509 c1_i_req_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3140_ net155 net154 net157 net156 _0890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_78_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3071_ _0836_ net470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4275__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4990__I net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6183__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _0403_ clknet_leaf_45_core_clock dmmu1.page_table\[10\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6761_ _0334_ clknet_leaf_36_core_clock dmmu0.page_table\[5\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5775__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3973_ _1631_ _1634_ _1635_ _1636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_53_Right_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7078__I net362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5712_ _2065_ _2743_ _2745_ net1098 _2751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_85_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6692_ _0265_ clknet_leaf_92_core_clock immu_1.high_addr_off\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5527__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5643_ _2711_ _0341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5574_ _2672_ _0311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold201 dmmu1.page_table\[9\]\[3\] net935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4525_ _1861_ _2033_ _2035_ dmmu1.page_table\[14\]\[6\] _2042_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold212 dmmu1.page_table\[7\]\[8\] net946 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold223 immu_1.page_table\[10\]\[3\] net957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5326__I net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold234 dmmu0.page_table\[4\]\[5\] net968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3274__C _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold245 dmmu0.page_table\[4\]\[6\] net979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4456_ _2000_ _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_40_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold256 dmmu0.page_table\[3\]\[0\] net990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold267 immu_1.page_table\[12\]\[10\] net1001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_62_Right_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold278 dmmu1.page_table\[6\]\[1\] net1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_leaf_103_core_clock_I clknet_4_2__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6711__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold289 dmmu1.page_table\[9\]\[0\] net1023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3407_ dmmu0.page_table\[4\]\[9\] dmmu0.page_table\[5\]\[9\] dmmu0.page_table\[6\]\[9\]
+ dmmu0.page_table\[7\]\[9\] _0871_ _0866_ _1148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7175_ net211 net639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3936__S1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4387_ _1839_ _1873_ _1909_ _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_42_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input245_I dcache_wb_adr[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6126_ _2989_ _0546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3338_ net151 dmmu1.long_off_reg\[1\] _1081_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6057_ _2794_ _2941_ _2943_ dmmu1.page_table\[2\]\[7\] _2951_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3269_ net1 _1014_ _1015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6861__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5008_ _2340_ _0077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6007__A2 _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4018__A1 _1654_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_71_Right_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5215__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5766__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4569__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6959_ _0532_ clknet_leaf_64_core_clock dmmu1.page_table\[1\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_53_core_clock_I clknet_4_15__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3872__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6241__CLK clknet_leaf_96_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Right_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4140__I net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6391__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output631_I net631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3552__I0 net138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4257__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5206__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5509__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4980__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3375__B _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6734__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4732__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4310_ _1770_ _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_10_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5290_ _2508_ _0191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4241_ _1867_ _0592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_1460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3299__A2 _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4040__S0 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_7_0_core_clock clknet_0_core_clock clknet_3_7_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4172_ _1811_ _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3123_ dmmu0.page_table\[12\]\[0\] dmmu0.page_table\[13\]\[0\] dmmu0.page_table\[14\]\[0\]
+ dmmu0.page_table\[15\]\[0\] _0872_ _0868_ _0873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_3054_ _0827_ net477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_2664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5748__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6813_ _0386_ clknet_leaf_44_core_clock dmmu1.page_table\[11\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_82_2675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_2686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6264__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3956_ immu_1.page_table\[4\]\[7\] immu_1.page_table\[5\]\[7\] immu_1.page_table\[6\]\[7\]
+ immu_1.page_table\[7\]\[7\] _1404_ _1540_ _1619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_46_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6744_ _0317_ clknet_leaf_69_core_clock dmmu1.page_table\[15\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_2096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3223__A2 _0961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6675_ _0248_ clknet_leaf_37_core_clock dmmu0.page_table\[2\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3887_ _1422_ _1546_ _1551_ _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_33_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5626_ _1796_ _2699_ _2701_ dmmu0.page_table\[5\]\[1\] _2703_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input195_I c1_sr_bus_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5557_ net95 _2646_ _2648_ dmmu0.page_table\[3\]\[12\] _2662_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_83_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input362_I ic1_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4508_ _2030_ _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_13_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _2623_ _0274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_1989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input56_I c0_o_mem_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4895__I _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4439_ _1815_ _1979_ _1982_ dmmu0.page_table\[0\]\[7\] _1990_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4487__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5684__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7158_ net172 net628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6109_ _1851_ _2975_ _2977_ dmmu1.page_table\[0\]\[3\] _2981_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7089_ net343 net496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5436__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_1290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5987__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6607__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3240__S _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4411__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6757__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output679_I net679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4714__A2 _2156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5911__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7181__I net400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3525__I0 net134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6287__CLK clknet_leaf_40_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4650__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3810_ _1405_ immu_1.page_table\[14\]\[2\] _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ _1819_ _2191_ _2193_ net984 _2203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_18 net397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_29 net261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3741_ immu_1.page_table\[0\]\[0\] immu_1.page_table\[1\]\[0\] immu_1.page_table\[2\]\[0\]
+ immu_1.page_table\[3\]\[0\] _1409_ _1410_ _1411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_27_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6460_ _0033_ clknet_leaf_102_core_clock dmmu0.page_table\[9\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6155__A1 _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3672_ _1345_ _1346_ _1347_ net680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_1470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5411_ _2578_ _0242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6391_ _0773_ clknet_leaf_80_core_clock immu_1.page_table\[10\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_1560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5342_ _2451_ _2536_ _2538_ dmmu0.page_table\[15\]\[1\] _2540_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_80_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5273_ net104 _2486_ _2488_ immu_0.page_table\[1\]\[9\] _2498_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_71_2354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4469__A1 _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4013__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4224_ _1854_ _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_23_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5130__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3141__A1 net151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4155_ net97 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_58_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3692__A2 net365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3106_ net50 net49 net52 net51 _0856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4086_ _1744_ _1712_ _1745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5969__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6091__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3037_ net388 _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_78_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input110_I c1_o_instr_long_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_2158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input208_I c1_sr_bus_data_o[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_2169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3995__S _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_2082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5197__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4988_ _2277_ _2317_ _2319_ net1079 _2327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_1835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_inner_713 c0_i_core_int_sreg[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_18_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinterconnect_inner_724 c1_i_core_int_sreg[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_6727_ _0300_ clknet_leaf_39_core_clock dmmu0.page_table\[3\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4944__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3939_ _1440_ _1602_ _1603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6170__I _3015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_Left_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_22_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_2069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6658_ _0231_ clknet_leaf_25_core_clock dmmu0.page_table\[11\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4157__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5609_ _2692_ _0326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6589_ _0162_ clknet_leaf_22_core_clock immu_0.page_table\[3\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3235__S _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput670 net670 inner_wb_adr[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput681 net681 inner_wb_adr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput692 net692 inner_wb_o_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3034__I _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4880__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3683__A2 net378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4632__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Left_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_1655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4935__A2 _2290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7176__I net389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput16 c0_o_mem_addr[12] net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput27 c0_o_mem_addr[8] net27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_68_1544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput38 c0_o_mem_data[3] net38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput49 c0_o_mem_high_addr[4] net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5360__A2 _2535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3653__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5112__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3674__A2 net376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6922__CLK clknet_leaf_64_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6073__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5960_ _2896_ _0473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4911_ _2277_ _2261_ _2263_ net943 _2278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5891_ _2682_ _2855_ _2857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_2011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4842_ _2234_ _0017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_2033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_16_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4773_ _2194_ _0797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4926__A2 _2137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3724_ _1385_ immu_0.page_table\[7\]\[0\] _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6512_ _0085_ clknet_leaf_6_core_clock immu_0.page_table\[10\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6302__CLK clknet_leaf_96_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_2541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3655_ _1332_ _1333_ _1334_ net676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6443_ _0016_ clknet_leaf_15_core_clock dmmu0.page_table\[10\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_2405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_73_2416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6374_ _0756_ clknet_leaf_73_core_clock immu_1.page_table\[11\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3586_ _1293_ net426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3362__A1 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5325_ _2528_ _0206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_1986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6452__CLK clknet_leaf_17_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input158_I c1_o_mem_long_mode vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5103__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5256_ _2489_ _0176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4207_ _1771_ _1840_ _1842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_3_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5187_ _2443_ _0153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3665__A2 net374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4862__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4138_ net82 net81 _1783_ _1784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_74_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input19_I c0_o_mem_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4069_ _1684_ _1727_ _1728_ _1729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4917__A2 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6119__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5342__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3353__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3656__A2 net372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6055__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4605__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5802__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6325__CLK clknet_leaf_70_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4908__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5419__I _2583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5581__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6475__CLK clknet_leaf_103_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3440_ net50 dmmu0.long_off_reg\[5\] _1180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3371_ dmmu0.page_table\[0\]\[8\] dmmu0.page_table\[1\]\[8\] dmmu0.page_table\[2\]\[8\]
+ dmmu0.page_table\[3\]\[8\] _0872_ _0941_ _1113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5110_ _2140_ _2397_ _2399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6090_ _2969_ _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_108_core_clock_I clknet_4_0__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5097__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5041_ _2271_ _2352_ _2354_ net1107 _2359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4993__I net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6992_ _0565_ clknet_leaf_94_core_clock dmmu1.long_off_reg\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_18_core_clock clknet_4_4__leaf_core_clock clknet_leaf_18_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5943_ _2851_ _2872_ _2874_ net774 _2886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_1796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5874_ _2794_ _2836_ _2838_ dmmu1.page_table\[8\]\[7\] _2846_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_2052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_2603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4825_ _1980_ _2223_ _2225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5021__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5329__I net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_58_core_clock_I clknet_4_14__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6818__CLK clknet_leaf_68_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4756_ _2183_ _0791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3583__A1 net228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4780__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3707_ net315 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4687_ _2141_ _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_43_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input275_I dcache_wb_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6426_ _0808_ clknet_leaf_110_core_clock immu_0.page_table\[13\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3638_ _1322_ net689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5324__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3335__A1 _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3335__B2 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3569_ net221 _1204_ _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6357_ _0739_ clknet_leaf_77_core_clock immu_1.page_table\[13\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5308_ _2519_ _0198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6288_ _0670_ clknet_leaf_13_core_clock dmmu0.page_table\[0\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput206 c1_sr_bus_data_o[6] net206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_57_core_clock clknet_4_14__leaf_core_clock clknet_leaf_57_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput217 dcache_mem_o_data[12] net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput228 dcache_mem_o_data[8] net228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput239 dcache_wb_adr[17] net239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5239_ _2478_ _0170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4835__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_110_core_clock_I clknet_4_0__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output494_I net494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6498__CLK clknet_leaf_32_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5563__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output661_I net661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_96_core_clock clknet_4_9__leaf_core_clock clknet_leaf_96_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5315__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3326__A1 net151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4523__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_60_core_clock_I clknet_4_14__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_2019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5079__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3629__A2 net271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold5 immu_1.page_table\[15\]\[4\] net739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_76_1621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5251__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Left_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_1248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4610_ _2095_ _0733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5590_ _2680_ _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_5_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3565__A1 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4541_ _1823_ _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_25_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4472_ _2009_ _0681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3317__A1 net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6211_ _0593_ clknet_leaf_80_core_clock immu_1.page_table\[9\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3423_ _0896_ _1163_ _1164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7191_ net395 net648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3868__A2 _1532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6142_ _2999_ _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_42_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3354_ dmmu0.page_table\[0\]\[7\] dmmu0.page_table\[1\]\[7\] dmmu0.page_table\[2\]\[7\]
+ dmmu0.page_table\[3\]\[7\] _0950_ _0952_ _1097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_29_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6073_ _2776_ _2958_ _2960_ net857 _2961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3285_ _0948_ _1027_ _1030_ _0940_ _1031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_77_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3176__S0 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5024_ _2348_ _0085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_1841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6019__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4293__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4228__I _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3132__I _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6975_ _0548_ clknet_leaf_105_core_clock mem_dcache_arb.select vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5242__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5926_ _2877_ _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6640__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5857_ _2835_ _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_14_1479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input392_I inner_wb_i_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4808_ _1806_ _2208_ _2210_ immu_0.page_table\[13\]\[4\] _2215_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5545__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5788_ _2103_ _2778_ _2780_ net1090 _2797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input86_I c0_sr_bus_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6790__CLK clknet_leaf_42_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4898__I _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4753__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4739_ _2171_ net76 _2172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_71_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6409_ _0791_ clknet_leaf_0_core_clock immu_0.page_table\[14\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3859__A2 _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4808__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5481__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output507_I net507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5784__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_1019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7184__I net403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6513__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3070_ net217 _0831_ _0836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_2016 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5224__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6760_ _0333_ clknet_leaf_48_core_clock dmmu0.page_table\[5\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5775__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3972_ _1631_ _1634_ net2 _1635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5711_ _2750_ _0370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3330__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6691_ _0264_ clknet_4_8__leaf_core_clock immu_1.high_addr_off\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5642_ _2529_ _2699_ _2701_ net787 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5527__A2 _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3836__B _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ _2065_ _2664_ _2666_ net949 _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold202 immu_1.page_table\[9\]\[5\] net936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4524_ _2041_ _0701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold213 dmmu0.page_table\[2\]\[6\] net947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold224 immu_0.page_table\[5\]\[3\] net958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold235 dmmu0.page_table\[2\]\[11\] net969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold246 immu_0.page_table\[8\]\[9\] net980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4455_ _1895_ _1998_ _2000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold257 dmmu0.page_table\[13\]\[10\] net991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold268 dmmu0.page_table\[12\]\[10\] net1002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold279 dmmu1.page_table\[0\]\[5\] net1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6193__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3406_ _1145_ _1146_ _0877_ _1147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7174_ net163 net638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4386_ _1955_ _0649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3337_ net151 dmmu1.long_off_reg\[1\] _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6125_ net199 _2974_ _2976_ dmmu1.page_table\[0\]\[11\] _2989_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_8_core_clock clknet_4_1__leaf_core_clock clknet_leaf_8_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input140_I c1_o_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input238_I dcache_wb_adr[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3268_ net53 _1014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6056_ _2950_ _0515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_1248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5007_ _2258_ _2337_ _2339_ immu_0.page_table\[10\]\[0\] _2340_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3199_ _0867_ _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_68_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5215__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5766__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6958_ _0531_ clknet_leaf_63_core_clock dmmu1.page_table\[1\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_104_core_clock clknet_4_2__leaf_core_clock clknet_leaf_104_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3321__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4974__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ _2847_ _2856_ _2858_ net946 _2867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6889_ _0462_ clknet_leaf_56_core_clock dmmu1.page_table\[6\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3872__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4726__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4421__I _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output457_I net457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5453__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3388__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5151__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3552__I1 net33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output624_I net624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6686__CLK clknet_leaf_92_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4257__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7179__I net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5206__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_2044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3768__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3312__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5509__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5390__B1 _2554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3940__A1 _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4240_ _1866_ _1841_ _1843_ immu_1.page_table\[9\]\[8\] _1867_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4040__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4171_ net101 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3122_ _0871_ _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3053_ net224 _0822_ _0827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_26_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6812_ _0385_ clknet_leaf_52_core_clock dmmu1.page_table\[11\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_82_2665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5748__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_2687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6743_ _0316_ clknet_leaf_42_core_clock dmmu1.page_table\[15\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4956__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3955_ immu_1.page_table\[0\]\[7\] immu_1.page_table\[1\]\[7\] immu_1.page_table\[2\]\[7\]
+ immu_1.page_table\[3\]\[7\] _1404_ _1540_ _1618_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_18_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_2097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6674_ _0247_ clknet_leaf_37_core_clock dmmu0.page_table\[2\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3886_ net107 _1549_ _1550_ _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6559__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5625_ _2702_ _0332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5337__I _2535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input188_I c1_sr_bus_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3285__C _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5556_ _2661_ _0304_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4507_ _1769_ _1837_ _2029_ _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_0_28_1968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5487_ _2463_ _2613_ _2615_ dmmu0.page_table\[4\]\[7\] _2623_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input355_I ic1_mem_data[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4438_ _1989_ _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4487__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5684__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input49_I c0_o_mem_high_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7157_ net171 net627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4369_ _1849_ _1942_ _1944_ immu_1.page_table\[4\]\[2\] _1947_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_67_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6108_ _2980_ _0537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7088_ net341 net494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5436__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6039_ _1891_ _1909_ _2030_ _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_9_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5987__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_46_1594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5372__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5911__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_2037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3922__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5124__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4650__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_19 net397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3740_ net367 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_12_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6155__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3671_ _1337_ net251 _1347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5410_ immu_0.high_addr_off\[5\] _1809_ _2572_ _2578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_11_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6851__CLK clknet_leaf_41_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6390_ _0772_ clknet_leaf_75_core_clock immu_1.page_table\[10\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3913__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4996__I net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5341_ _2539_ _0211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_75_2480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5272_ _2497_ _0184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_71_2355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4013__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4469__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4223_ net204 _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3141__A2 net150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4154_ _1798_ _0574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5418__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3105_ _0855_ net519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6231__CLK clknet_leaf_85_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4085_ net11 immu_0.high_addr_off\[6\] _1744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5969__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6091__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3036_ _0812_ _0814_ _0815_ net602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_84_2749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4236__I _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_2037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input103_I c0_sr_bus_data_o[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6381__CLK clknet_leaf_73_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4987_ _2326_ _0070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_1983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinterconnect_inner_714 c0_i_core_int_sreg[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_18_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6726_ _0299_ clknet_leaf_40_core_clock dmmu0.page_table\[3\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3938_ immu_1.page_table\[0\]\[6\] immu_1.page_table\[1\]\[6\] immu_1.page_table\[2\]\[6\]
+ immu_1.page_table\[3\]\[6\] _1474_ _1433_ _1602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_74_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinterconnect_inner_725 c1_i_core_int_sreg[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_22_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6657_ _0230_ clknet_leaf_16_core_clock dmmu0.page_table\[11\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3869_ inner_wb_arbiter.o_sel_sig _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_2_1093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4157__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5608_ _2463_ _2681_ _2684_ net1029 _2692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5354__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6588_ _0161_ clknet_leaf_17_core_clock immu_0.page_table\[3\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3904__A1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5539_ _2455_ _2647_ _2649_ net952 _2653_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput660 net660 inner_wb_adr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_2081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput671 net671 inner_wb_adr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_54_1841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput682 net682 inner_wb_adr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput693 net693 inner_wb_o_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_65_core_clock_I clknet_4_15__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4880__A2 _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5530__I _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6724__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6874__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput17 c0_o_mem_addr[13] net17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 c0_o_mem_addr[9] net28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_68_1556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput39 c0_o_mem_data[4] net39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_1767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5648__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6254__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3754__S0 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5820__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4910_ _1814_ _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_34_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5890_ _2855_ _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_73_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_2012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _1815_ _2224_ _2226_ net932 _2234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_2023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4387__A1 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4772_ _1777_ _2191_ _2193_ net995 _2194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_16_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4926__A3 _2286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6511_ _0084_ clknet_leaf_5_core_clock immu_0.page_table\[10\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3723_ _1372_ _1388_ _1389_ _1392_ _1367_ _1393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XTAP_TAPCELL_ROW_77_2520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6442_ _0015_ clknet_leaf_24_core_clock dmmu0.page_table\[10\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3654_ _1306_ net247 _1334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_2406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5887__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_2417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6373_ _0755_ clknet_leaf_96_core_clock immu_1.page_table\[11\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3585_ net229 _1219_ _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_60_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5324_ _2527_ _2516_ _2518_ dmmu0.page_table\[12\]\[8\] _2528_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3993__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_47_core_clock clknet_4_13__leaf_core_clock clknet_leaf_47_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5255_ _1776_ _2486_ _2488_ immu_0.page_table\[1\]\[0\] _2489_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4311__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4206_ _1840_ _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_3_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5186_ _2332_ _2429_ _2431_ net1068 _2443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_3_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4862__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4137_ net80 net79 net78 net77 _1783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA_input220_I dcache_mem_o_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input318_I ic0_wb_adr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4068_ net115 immu_1.high_addr_off\[5\] _1728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_39_1179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5662__I1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6897__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5414__I1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_43_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5575__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6709_ _0282_ clknet_leaf_33_core_clock dmmu0.page_table\[13\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3976__I1 _1638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6119__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_86_core_clock clknet_4_10__leaf_core_clock clknet_leaf_86_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5327__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6277__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput490 net490 c1_i_req_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6055__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5802__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7187__I net391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3041__A1 net559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3370_ _1110_ _1111_ _0938_ _1112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3975__S0 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5097__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5040_ _2358_ _0091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_2800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6991_ _0564_ clknet_leaf_94_core_clock dmmu1.long_off_reg\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_1622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5942_ _2885_ _0466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5873_ _2845_ _0437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3280__A1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4824_ _2223_ _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_12_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_2075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5021__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4755_ _1809_ _2175_ _2177_ immu_0.page_table\[14\]\[5\] _2183_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5309__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4780__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3583__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3706_ immu_0.page_table\[8\]\[0\] immu_0.page_table\[9\]\[0\] immu_0.page_table\[10\]\[0\]
+ immu_0.page_table\[11\]\[0\] _1370_ _1372_ _1376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_44_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4686_ _2140_ _2138_ _2141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6425_ _0807_ clknet_leaf_107_core_clock immu_0.page_table\[12\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3637_ _0812_ net260 _1322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input170_I c1_o_req_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input268_I dcache_wb_o_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3335__A2 _1076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6356_ _0738_ clknet_leaf_63_core_clock immu_1.page_table\[13\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3568_ _1284_ net411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5307_ _2444_ _2516_ _2518_ net925 _2519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6287_ _0669_ clknet_leaf_40_core_clock dmmu0.page_table\[0\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3499_ dmmu0.page_table\[0\]\[12\] dmmu0.page_table\[1\]\[12\] dmmu0.page_table\[2\]\[12\]
+ dmmu0.page_table\[3\]\[12\] _0863_ _0866_ _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xinput207 c1_sr_bus_data_o[7] net207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput218 dcache_mem_o_data[13] net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput229 dcache_mem_o_data[9] net229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5238_ _2459_ _2470_ _2472_ immu_0.page_table\[2\]\[5\] _2478_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input31_I c0_o_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4835__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5169_ _2434_ _0144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6037__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4599__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output487_I net487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4523__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4523__B2 dmmu1.page_table\[14\]\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5720__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4287__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold6 dmmu0.page_table\[7\]\[2\] net740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_76_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6442__CLK clknet_leaf_24_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5539__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5003__A2 _2222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_2073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_2084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3565__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ _2050_ _0708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6592__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4471_ _1863_ _1999_ _2001_ immu_1.page_table\[1\]\[7\] _2009_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_42_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6210_ _0592_ clknet_leaf_81_core_clock immu_1.page_table\[9\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3422_ dmmu1.page_table\[4\]\[9\] dmmu1.page_table\[5\]\[9\] dmmu1.page_table\[6\]\[9\]
+ dmmu1.page_table\[7\]\[9\] _0886_ _0900_ _1163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_42_2046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7190_ net394 net647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6141_ _1826_ _1839_ _1892_ _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3353_ _0940_ _1095_ _1096_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6072_ _2959_ _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3284_ _0882_ _1028_ _1029_ _0948_ _1030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_20_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5023_ _2328_ _2337_ _2339_ net1106 _2348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3176__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6019__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5778__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6974_ _0547_ clknet_leaf_64_core_clock dmmu1.page_table\[0\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_2115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5242__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5925_ _2782_ _2873_ _2875_ net1012 _2877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3253__A1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5856_ _1826_ _1892_ _2031_ _2835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_75_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_3_Right_3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4807_ _2214_ _0002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6935__CLK clknet_leaf_64_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5787_ _2796_ _0400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_1171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4753__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input385_I inner_embed_mode vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4738_ net83 _2171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input79_I c0_sr_bus_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4669_ _2130_ _0757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6408_ _0790_ clknet_leaf_112_core_clock immu_0.page_table\[14\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4505__A1 net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5702__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6339_ _0721_ clknet_leaf_76_core_clock immu_1.page_table\[14\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6315__CLK clknet_leaf_70_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4269__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4808__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4419__I _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5481__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3492__A1 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3492__B2 _1119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6465__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5769__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4441__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3198__C _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4044__I0 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5941__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6808__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_2006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3322__I2 dmmu1.page_table\[14\]\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3483__A1 _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6958__CLK clknet_leaf_63_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3971_ _1632_ _1633_ _1634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5710_ _2063_ _2743_ _2745_ dmmu1.page_table\[12\]\[4\] _2750_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6690_ _0263_ clknet_leaf_92_core_clock immu_1.high_addr_off\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3330__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5641_ _2710_ _0340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5572_ _2671_ _0310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4523_ _1858_ _2033_ _2035_ dmmu1.page_table\[14\]\[5\] _2041_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold203 dmmu0.page_table\[15\]\[10\] net937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold214 immu_1.page_table\[4\]\[5\] net948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold225 dmmu1.page_table\[12\]\[3\] net959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4454_ _1998_ _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6338__CLK clknet_leaf_63_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold236 immu_0.page_table\[6\]\[9\] net970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold247 dmmu1.page_table\[0\]\[0\] net981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4499__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold258 dmmu0.page_table\[2\]\[5\] net992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold269 dmmu1.page_table\[5\]\[9\] net1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3405_ dmmu0.page_table\[8\]\[9\] dmmu0.page_table\[9\]\[9\] dmmu0.page_table\[10\]\[9\]
+ dmmu0.page_table\[11\]\[9\] _0871_ _0866_ _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7173_ net180 net637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4385_ _1870_ _1941_ _1943_ immu_1.page_table\[4\]\[10\] _1955_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3171__B1 _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6124_ _2988_ _0545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3336_ _1071_ _1079_ net526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__4239__I net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6488__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6055_ _2792_ _2941_ _2943_ net802 _2950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3267_ net124 _0933_ _0989_ _1012_ _0841_ _1013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__5999__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input133_I c1_o_mem_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5006_ _2338_ _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3474__A1 _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3198_ _0879_ _0939_ _0946_ _0883_ _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_7_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input300_I ic0_mem_data[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5215__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_2081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6957_ _0530_ clknet_leaf_62_core_clock dmmu1.page_table\[1\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4974__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3321__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5908_ _2866_ _0451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6888_ _0461_ clknet_leaf_59_core_clock dmmu1.page_table\[6\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5839_ _2826_ _0422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_1919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4726__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Left_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5151__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3388__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3254__S _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_24_Left_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5206__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3217__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3312__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_72_core_clock_I clknet_4_9__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4193__A2 net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5390__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6630__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4170_ _1810_ _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3121_ _0863_ _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3052_ _0826_ net476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6780__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput390 inner_wb_i_dat[10] net390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_37_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6811_ _0384_ clknet_leaf_50_core_clock dmmu1.page_table\[11\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_2666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4405__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_2688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6742_ _0315_ clknet_leaf_42_core_clock dmmu1.page_table\[15\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4956__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3954_ net113 immu_1.high_addr_off\[3\] _1616_ _1617_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_19_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_2098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6673_ _0246_ clknet_leaf_41_core_clock dmmu0.page_table\[2\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3885_ _1547_ _1548_ _1550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5624_ _1776_ _2699_ _2701_ dmmu0.page_table\[5\]\[0\] _2702_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_27_972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4708__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5905__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5555_ net94 _2646_ _2648_ dmmu0.page_table\[3\]\[11\] _2661_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3138__I _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4506_ _1830_ net196 _1831_ _1832_ _2029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5486_ _2622_ _0273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4437_ _1812_ _1979_ _1982_ net904 _1989_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input250_I dcache_wb_adr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input348_I ic1_mem_data[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5684__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7156_ net164 net620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4368_ _1946_ _0640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6107_ _1848_ _2975_ _2977_ net1100 _2980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3319_ _1052_ _1063_ net525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7087_ net340 net493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4299_ _1863_ _1894_ _1897_ immu_1.page_table\[0\]\[7\] _1905_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_52_1780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5436__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6038_ _2939_ _0508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3447__A1 net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4644__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_2007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6149__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3249__S _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5372__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6653__CLK clknet_leaf_17_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_1473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3922__A2 _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5124__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3438__A1 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3670_ _0814_ net321 _1326_ _1346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_1595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5340_ _2444_ _2536_ _2538_ dmmu0.page_table\[15\]\[0\] _2539_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_51_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3913__A2 net239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_2470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_2481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5271_ net103 _2486_ _2488_ immu_0.page_table\[1\]\[8\] _2497_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xclkbuf_leaf_37_core_clock clknet_4_7__leaf_core_clock clknet_leaf_37_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_71_2334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4222_ _1853_ _0587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3677__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3141__A3 net153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4153_ _1797_ _1792_ _1794_ net751 _1798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5418__A2 _2581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3104_ net119 net14 _0850_ _0855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_1306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4084_ _1306_ _1725_ _1742_ _1743_ net674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__3429__A1 _1154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6091__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_2274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3035_ net387 _0815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_TAPCELL_ROW_69_2296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_1096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4986_ _2275_ _2317_ _2319_ net1016 _2326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5051__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3937_ _1434_ _1600_ _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6725_ _0298_ clknet_leaf_38_core_clock dmmu0.page_table\[3\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinterconnect_inner_715 c0_i_core_int_sreg[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_19_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinterconnect_inner_726 c1_i_core_int_sreg[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_73_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6676__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input298_I ic0_mem_data[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6656_ _0229_ clknet_leaf_25_core_clock dmmu0.page_table\[11\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3868_ _1382_ _1532_ _1533_ net2 _1422_ _1534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xclkbuf_leaf_76_core_clock clknet_4_11__leaf_core_clock clknet_leaf_76_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_12__f_core_clock clknet_3_6_0_core_clock clknet_4_12__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_27_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _2691_ _0325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5354__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4157__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ _0160_ clknet_leaf_18_core_clock immu_0.page_table\[3\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3799_ _1375_ _1381_ _1466_ _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_28_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5538_ _2652_ _0295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input61_I c0_o_req_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5469_ _1976_ _2428_ _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xoutput650 net650 ic1_wb_i_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput661 net661 inner_wb_adr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput672 net672 inner_wb_adr[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput683 net683 inner_wb_adr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput694 net694 inner_wb_o_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7139_ net211 net601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4617__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_48_1646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5459__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 c0_o_mem_addr[14] net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput29 c0_o_mem_data[0] net29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_1508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5648__A2 _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3203__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3659__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3754__S1 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6549__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6073__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4084__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3831__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4840_ _2233_ _0016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_60_2013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_2024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3397__B _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4387__A2 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4771_ _2192_ _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_16_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6510_ _0083_ clknet_leaf_6_core_clock immu_0.page_table\[10\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3722_ _1385_ immu_0.page_table\[3\]\[0\] _1391_ _1392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_82_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_2521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6441_ _0014_ clknet_leaf_38_core_clock dmmu0.page_table\[10\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_2543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3653_ _0814_ net317 _1326_ _1333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6372_ _0754_ clknet_leaf_75_core_clock immu_1.page_table\[11\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3584_ _1292_ net425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_1321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_2066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3898__A1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5323_ net103 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3993__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5254_ _2487_ _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4847__B1 _2225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4205_ _1829_ _1839_ _1840_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5185_ _2442_ _0152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_3_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4136_ net91 _1782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_79_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4067_ net115 immu_1.high_addr_off\[5\] _1727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3151__I _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input213_I dcache_mem_exception vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5575__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4969_ _2315_ _0063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_1167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6708_ _0281_ clknet_leaf_29_core_clock dmmu0.page_table\[13\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5327__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6639_ _0212_ clknet_leaf_28_core_clock dmmu0.page_table\[15\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3527__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3889__A1 net6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput480 net480 c1_i_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput491 net491 c1_i_req_data[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_output432_I net432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6055__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3061__I _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4066__A1 net116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6841__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5263__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5802__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3813__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5015__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_11_core_clock_I clknet_4_3__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6991__CLK clknet_leaf_94_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4106__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6221__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3424__S0 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3975__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5652__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6371__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4829__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3680__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_2200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4057__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6990_ _0563_ clknet_leaf_104_core_clock inner_wb_arbiter.o_sel_sig vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_36_1309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3104__I0 net119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5941_ _2849_ _2873_ _2875_ net876 _2885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5872_ _2792_ _2836_ _2838_ net1062 _2845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _1977_ _2222_ _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_29_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5557__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4754_ _2182_ _0790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5309__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3705_ _1366_ _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_71_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4780__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4685_ _1770_ _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6424_ _0806_ clknet_leaf_0_core_clock immu_0.page_table\[12\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3636_ _1321_ net688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6714__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6355_ _0737_ clknet_leaf_76_core_clock immu_1.page_table\[13\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3567_ net214 _1204_ _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3146__I net122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input163_I c1_o_req_active vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5306_ _2517_ _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_12_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6286_ _0668_ clknet_leaf_40_core_clock dmmu0.page_table\[0\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3498_ net52 dmmu0.long_off_reg\[7\] _1235_ _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
Xinput208 c1_sr_bus_data_o[8] net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5237_ _2477_ _0169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput219 dcache_mem_o_data[14] net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input330_I ic1_mem_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_core_clock_I core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5168_ _2265_ _2430_ _2432_ immu_0.page_table\[4\]\[1\] _2434_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input24_I c0_o_mem_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6037__A2 _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4119_ _1772_ net462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4048__A1 net11 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5099_ _2277_ _2382_ _2384_ immu_0.page_table\[7\]\[7\] _2392_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5796__A1 _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_2_core_clock_I clknet_4_1__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6244__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_77_core_clock_I clknet_4_11__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3484__C _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4523__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5720__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4287__A1 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold7 immu_1.page_table\[10\]\[8\] net741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_57_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__A1 net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5236__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_2065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3893__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5539__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6737__CLK clknet_leaf_46_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4470_ _2008_ _0680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3421_ _1160_ _1161_ _0906_ _1162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_81_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6887__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6140_ _2998_ _0551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3352_ dmmu0.page_table\[4\]\[7\] dmmu0.page_table\[5\]\[7\] dmmu0.page_table\[6\]\[7\]
+ dmmu0.page_table\[7\]\[7\] _0882_ _0948_ _1095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_21_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6071_ _1770_ _2957_ _2959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3283_ _0865_ dmmu0.page_table\[8\]\[4\] _1029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5475__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5022_ _2347_ _0084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6019__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5778__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6973_ _0546_ clknet_leaf_65_core_clock dmmu1.page_table\[0\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6267__CLK clknet_leaf_89_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5924_ _2876_ _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5855_ _2834_ _0430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4806_ _1803_ _2208_ _2210_ net1059 _2214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5786_ _2101_ _2778_ _2780_ net986 _2796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4737_ _2170_ _0785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4753__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input280_I ic0_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input378_I ic1_wb_adr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4668_ _2063_ _2123_ _2125_ immu_1.page_table\[11\]\[4\] _2130_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6407_ _0789_ clknet_leaf_108_core_clock immu_0.page_table\[14\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3619_ _1308_ net266 _1313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4505__A2 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5702__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4599_ _1870_ _2074_ _2076_ net907 _2088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4061__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6338_ _0720_ clknet_leaf_63_core_clock immu_1.page_table\[14\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6269_ _0651_ clknet_leaf_87_core_clock immu_1.page_table\[6\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4269__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3540__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5769__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4441__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output597_I net597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5467__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_2014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5941__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Right_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5209__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4680__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3970_ net8 immu_0.high_addr_off\[3\] _1633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5640_ _2527_ _2699_ _2701_ net996 _2710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_2114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5571_ _2063_ _2664_ _2666_ net870 _2671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4522_ _2040_ _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold204 dmmu1.page_table\[8\]\[12\] net938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_48_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold215 dmmu1.page_table\[15\]\[5\] net949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold226 dmmu0.page_table\[13\]\[3\] net960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4453_ _1828_ _1838_ _1891_ _1998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
Xhold237 dmmu1.page_table\[4\]\[1\] net971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4499__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4043__S0 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold248 immu_1.page_table\[12\]\[7\] net982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3546__I0 net135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold259 immu_1.page_table\[14\]\[9\] net993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3404_ dmmu0.page_table\[12\]\[9\] dmmu0.page_table\[13\]\[9\] dmmu0.page_table\[14\]\[9\]
+ dmmu0.page_table\[15\]\[9\] _0871_ _0867_ _1145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7172_ net109 net636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4384_ _1954_ _0648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3171__A1 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6123_ _2851_ _2974_ _2976_ dmmu1.page_table\[0\]\[10\] _2988_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3335_ _0862_ _1076_ _1078_ _0860_ _0884_ _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_42_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6054_ _2949_ _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_31_Right_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5999__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3266_ _0915_ _0994_ _0999_ _1004_ _1011_ _1012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_77_1228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5005_ _2140_ _2336_ _2338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3197_ _0943_ _0945_ _0879_ _0946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__3474__A2 _1212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input126_I c1_o_mem_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6956_ _0529_ clknet_leaf_57_core_clock dmmu1.page_table\[1\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ _2794_ _2856_ _2858_ net1046 _2866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4974__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6887_ _0460_ clknet_leaf_55_core_clock dmmu1.page_table\[6\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Right_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5838_ _1805_ _2819_ _2821_ dmmu0.page_table\[1\]\[4\] _2826_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input91_I c0_sr_bus_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5769_ _2784_ _2778_ _2780_ dmmu1.page_table\[10\]\[2\] _2785_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3785__I0 net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5151__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6432__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output512_I net512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4662__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6582__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3217__A2 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4414__A1 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1946 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6167__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5390__A2 _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4025__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_27_core_clock clknet_4_5__leaf_core_clock clknet_leaf_27_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5678__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5660__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3120_ dmmu0.page_table\[0\]\[0\] dmmu0.page_table\[1\]\[0\] dmmu0.page_table\[2\]\[0\]
+ dmmu0.page_table\[3\]\[0\] _0865_ _0868_ _0870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6925__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3051_ net223 _0822_ _0826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput380 ic1_wb_sel[0] net380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput391 inner_wb_i_dat[11] net391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5850__B1 _2820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6810_ _0383_ clknet_leaf_52_core_clock dmmu1.page_table\[11\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4405__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5602__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_2678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_2689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6741_ _0314_ clknet_leaf_45_core_clock dmmu1.page_table\[15\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3953_ _1613_ _1615_ _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4956__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_2099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3884_ _1547_ _1548_ _1549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6672_ _0245_ clknet_leaf_38_core_clock dmmu0.page_table\[2\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6305__CLK clknet_leaf_89_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_66_core_clock clknet_4_12__leaf_core_clock clknet_leaf_66_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4169__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5905__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5623_ _2700_ _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_73_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5554_ _2660_ _0303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4505_ net190 net189 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_44_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5485_ _2461_ _2613_ _2615_ net979 _2622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6455__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4436_ _1988_ _0666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6181__I1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3144__A1 net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4341__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4367_ _1846_ _1942_ _1944_ immu_1.page_table\[4\]\[1\] _1946_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7155_ net395 net610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input243_I dcache_wb_adr[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6106_ _2979_ _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3318_ _0862_ _1061_ _1062_ _0860_ _0884_ _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7086_ net339 net492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4298_ _1904_ _0612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_52_1770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6037_ net200 _2923_ _2925_ net807 _2939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_52_1792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3249_ dmmu1.page_table\[2\]\[4\] dmmu1.page_table\[3\]\[4\] _0908_ _0995_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_1913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4644__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6939_ _0512_ clknet_leaf_54_core_clock dmmu1.page_table\[2\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4713__I _2156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6149__A1 _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_16_core_clock_I clknet_4_6__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5372__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3383__A1 net152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output462_I net462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_2039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5124__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3135__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6948__CLK clknet_leaf_64_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6085__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5832__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6328__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4399__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_1__f_core_clock clknet_3_0_0_core_clock clknet_4_1__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_3_1530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6478__CLK clknet_leaf_32_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5899__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3374__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4571__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3175__S _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5270_ _2496_ _0183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4323__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4221_ _1852_ _1841_ _1843_ immu_1.page_table\[9\]\[3\] _1853_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_27_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3677__A2 net252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4152_ _1796_ _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3141__A4 net152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_2019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3103_ _0854_ net541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4083_ _1535_ net245 _1743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3702__I _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3034_ _0813_ _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_84_2729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_Left_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4929__A2 _2240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4985_ _2325_ _0069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5051__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6724_ _0297_ clknet_leaf_38_core_clock dmmu0.page_table\[3\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3936_ immu_1.page_table\[4\]\[6\] immu_1.page_table\[5\]\[6\] immu_1.page_table\[6\]\[6\]
+ immu_1.page_table\[7\]\[6\] _1474_ _1433_ _1600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_50_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_inner_716 c0_i_core_int_sreg[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_clkbuf_leaf_7_core_clock_I clknet_4_1__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_inner_727 c1_i_core_int_sreg[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_18_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6655_ _0228_ clknet_leaf_31_core_clock dmmu0.page_table\[11\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3867_ net5 immu_0.high_addr_off\[0\] _1533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3149__I _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input193_I c1_sr_bus_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5606_ _2461_ _2681_ _2684_ net771 _2691_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5354__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6586_ _0159_ clknet_leaf_24_core_clock immu_0.page_table\[3\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3798_ _1372_ _1461_ _1465_ _1377_ _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_14_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3365__A1 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5537_ _2453_ _2647_ _2649_ net833 _2652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3085__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input360_I ic1_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Left_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput640 net640 ic1_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5468_ _2611_ _0266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input54_I c0_o_mem_req vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput651 net651 ic1_wb_i_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput662 net662 inner_wb_adr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput673 net673 inner_wb_adr[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4419_ _1976_ _1977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput684 net684 inner_wb_cyc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput695 net695 inner_wb_o_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5399_ _2571_ _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_22_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_1707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7138_ net58 net600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7069_ net331 net484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4617__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5814__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_61_Left_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_1885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_48_1658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3768__B net705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 c0_o_mem_addr[15] net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_21_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_70_Left_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6770__CLK clknet_leaf_42_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3203__S1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3659__A2 net248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4856__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_84_core_clock_I clknet_4_10__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4084__A2 _1725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_2150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5033__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_2014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4387__A3 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4770_ _2140_ _2190_ _2192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_16_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3595__A1 net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3721_ _1390_ _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_71_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_2050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_2522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6440_ _0013_ clknet_leaf_31_core_clock dmmu0.page_table\[10\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_2533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3652_ _1302_ net371 _1332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_11__f_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3347__A1 _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_2408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3583_ net228 _1219_ _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6371_ _0753_ clknet_leaf_79_core_clock immu_1.page_table\[11\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_2419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5322_ _2526_ _0205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5253_ _1895_ _2485_ _2487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4847__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4204_ _1838_ _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5184_ _2330_ _2430_ _2432_ net961 _2442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6049__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4135_ _1779_ _1780_ _1781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_3_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4066_ net116 immu_1.high_addr_off\[6\] _1726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_39_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6643__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input206_I c1_sr_bus_data_o[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4968_ _1996_ _2298_ _2301_ net1065 _2315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5575__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6707_ _0280_ clknet_leaf_29_core_clock dmmu0.page_table\[13\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3130__S0 _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6793__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3919_ immu_0.page_table\[4\]\[6\] immu_0.page_table\[5\]\[6\] immu_0.page_table\[6\]\[6\]
+ immu_0.page_table\[7\]\[6\] _1424_ _1455_ _1583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_47_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4899_ _2269_ _2261_ _2263_ net804 _2270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6638_ _0211_ clknet_leaf_28_core_clock dmmu0.page_table\[15\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5327__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3338__A1 net151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6569_ _0142_ clknet_leaf_9_core_clock immu_0.page_table\[5\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_56_1905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput470 net470 c1_i_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput481 net481 c1_i_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput492 net492 c1_i_req_data[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3510__A1 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5263__A1 _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5015__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_69_Right_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3577__A1 net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_2018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4901__I _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3424__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_78_Right_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4829__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3188__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6666__CLK clknet_leaf_109_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_2802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_2201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_2212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3104__I1 net14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5940_ _2884_ _0465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_1646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5871_ _2844_ _0436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_1411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4822_ _1779_ _2172_ _2222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_34_1067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5557__A2 _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_1490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4016__C _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_2077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4753_ _1806_ _2175_ _2177_ immu_0.page_table\[14\]\[4\] _2182_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3704_ _1368_ _1373_ _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5309__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4684_ _2138_ _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_47_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6423_ _0805_ clknet_leaf_112_core_clock immu_0.page_table\[12\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4517__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3635_ _0812_ net259 _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_24_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6196__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6354_ _0736_ clknet_leaf_76_core_clock immu_1.page_table\[13\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3566_ _1283_ net410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_1715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5305_ _2300_ _2515_ _2517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_41_1016 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3497_ _1229_ _1233_ _1234_ _1235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6285_ _0667_ clknet_leaf_41_core_clock dmmu0.page_table\[0\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input156_I c1_o_mem_high_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput209 c1_sr_bus_data_o[9] net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_23_1450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5236_ _2457_ _2470_ _2472_ immu_0.page_table\[2\]\[4\] _2477_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5493__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5167_ _2433_ _0143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3162__I net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input323_I ic0_wb_adr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4118_ icore_sregs.c1_disable net384 _1772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5098_ _2391_ _0116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input17_I c0_o_mem_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4049_ net10 immu_0.high_addr_off\[5\] _1709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_78_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5796__A2 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3538__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6539__CLK clknet_leaf_6_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5720__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output542_I net542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6689__CLK clknet_leaf_91_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4287__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4168__I _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold8 dmmu1.page_table\[11\]\[8\] net742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5236__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3098__I0 net131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3798__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3342__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4117__B _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3893__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5539__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4747__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3970__A1 net8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_2015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3420_ dmmu1.page_table\[8\]\[9\] dmmu1.page_table\[9\]\[9\] dmmu1.page_table\[10\]\[9\]
+ dmmu1.page_table\[11\]\[9\] _0887_ _0900_ _1161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5172__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3722__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_2059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3351_ net106 net158 _0884_ _1093_ _1094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_1_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6070_ _2957_ _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3282_ dmmu0.page_table\[9\]\[4\] _1028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5475__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input9_I c0_o_instr_long_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5021_ _2277_ _2337_ _2339_ net773 _2347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3089__I0 net127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3710__I net3 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6972_ _0545_ clknet_leaf_64_core_clock dmmu1.page_table\[0\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5778__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5923_ _2776_ _2873_ _2875_ net839 _2876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4986__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5854_ net95 _2818_ _2820_ dmmu0.page_table\[1\]\[12\] _2834_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4805_ _2213_ _0001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5785_ _2795_ _0399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4541__I _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4736_ _1821_ _2156_ _2158_ net911 _2170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3961__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4667_ _2129_ _0756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3157__I _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input273_I dcache_wb_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6406_ _0788_ clknet_leaf_1_core_clock immu_0.page_table\[14\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6831__CLK clknet_leaf_68_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3618_ _1312_ net694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5702__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4598_ _2087_ _0729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4061__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6337_ _0719_ clknet_leaf_71_core_clock immu_1.page_table\[15\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3549_ _1274_ net545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3093__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6268_ _0650_ clknet_leaf_84_core_clock immu_1.page_table\[6\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4269__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6981__CLK clknet_leaf_96_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5219_ _2330_ _2447_ _2449_ net845 _2466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_2033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6199_ _0581_ clknet_leaf_6_core_clock immu_0.page_table\[11\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6211__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3324__S0 _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4441__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6361__CLK clknet_leaf_63_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output492_I net492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4044__I2 _1703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5941__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_1694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_17_core_clock clknet_4_5__leaf_core_clock clknet_leaf_17_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_31_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_1672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3704__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Left_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_1380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_23_core_clock_I clknet_4_4__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_2019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5209__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3530__I _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6704__CLK clknet_leaf_99_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5658__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_2104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_56_core_clock clknet_4_14__leaf_core_clock clknet_leaf_56_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_31_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6854__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5570_ _2670_ _0309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4521_ _1855_ _2033_ _2035_ dmmu1.page_table\[14\]\[4\] _2040_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold205 immu_1.page_table\[11\]\[3\] net939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_79_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5145__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4452_ _1997_ _0673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold216 dmmu1.page_table\[15\]\[2\] net950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold227 immu_0.page_table\[4\]\[9\] net961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold238 dmmu1.page_table\[13\]\[11\] net972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4499__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold249 immu_1.page_table\[12\]\[8\] net983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4043__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5696__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3546__I1 net30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3403_ _1119_ _1143_ _1144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_1723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7171_ net170 net626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4383_ _1868_ _1942_ _1944_ immu_1.page_table\[4\]\[9\] _1954_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_21_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3705__I _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3171__A2 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6122_ _2987_ _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3334_ net46 dmmu0.long_off_reg\[1\] _1077_ _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__5448__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6234__CLK clknet_leaf_96_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6053_ _2790_ _2941_ _2943_ net827 _2949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3265_ _0907_ _1007_ _1010_ _0912_ _1011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__5999__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4120__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5004_ _2336_ _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_56_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3196_ _0938_ _0944_ _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_95_core_clock clknet_4_8__leaf_core_clock clknet_leaf_95_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_1527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6384__CLK clknet_leaf_97_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_2059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input119_I c1_o_mem_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6955_ _0528_ clknet_leaf_58_core_clock dmmu1.page_table\[1\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5620__A1 _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4423__A2 _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5906_ _2865_ _0450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6886_ _0459_ clknet_leaf_51_core_clock dmmu1.page_table\[6\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_9__f_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5837_ _2825_ _0421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5367__I _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input390_I inner_wb_i_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5384__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5768_ _1848_ _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input84_I c0_sr_bus_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3934__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4719_ _2161_ _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3785__I1 _1453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5699_ _2742_ _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_60_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_2092 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_2076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6727__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4662__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output505_I net505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_89_core_clock_I clknet_4_8__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4414__A2 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_2085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6877__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6167__A2 net255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5277__I _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3925__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5678__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4025__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3050_ _0825_ net475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4102__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput370 ic1_wb_adr[1] net370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput381 ic1_wb_sel[1] net381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5850__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput392 inner_wb_i_dat[12] net392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_19_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4405__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5453__I1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_2679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6740_ _0313_ clknet_leaf_44_core_clock dmmu1.page_table\[15\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3952_ _1606_ _1549_ _1614_ _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6671_ _0244_ clknet_leaf_107_core_clock immu_0.high_addr_off\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3883_ net111 immu_1.high_addr_off\[1\] _1548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4169__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5622_ _2682_ _2698_ _2700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3216__I0 _0962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5905__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3916__A1 net6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5553_ _2531_ _2646_ _2648_ dmmu0.page_table\[3\]\[10\] _2660_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_91_core_clock_I clknet_4_8__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4504_ _2027_ _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5118__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5484_ _2621_ _0272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4435_ _1809_ _1979_ _1982_ net882 _1988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4341__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7154_ net394 net609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4366_ _1945_ _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6105_ _1845_ _2975_ _2977_ net902 _2979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3317_ net45 dmmu0.long_off_reg\[0\] _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7085_ net338 net491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4297_ _1860_ _1894_ _1897_ immu_1.page_table\[0\]\[6\] _1904_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_input236_I dcache_wb_adr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _2938_ _0507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_52_1793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3248_ _0931_ _0990_ _0993_ _0906_ _0994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4644__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3179_ _0907_ _0927_ _0928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input403_I inner_wb_i_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6938_ _0511_ clknet_leaf_53_core_clock dmmu1.page_table\[2\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6149__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6869_ _0442_ clknet_leaf_66_core_clock dmmu1.page_table\[8\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_46_1597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3546__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3135__A2 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output622_I net622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5560__I _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3281__S _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6085__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3518__S0 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4176__I _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3080__I _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4399__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4904__I _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5596__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_7_core_clock clknet_4_1__leaf_core_clock clknet_leaf_7_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5348__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5899__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4571__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_75_2461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_2483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4220_ _1851_ _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4323__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_2358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_103_core_clock clknet_4_2__leaf_core_clock clknet_leaf_103_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4874__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4151_ net96 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_2058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5470__I _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3102_ net133 net28 _0850_ _0854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4082_ _1422_ _1732_ _1741_ _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_39_1308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3033_ icache_arbiter.o_sel_sig _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_69_2276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5587__B1 _2665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4984_ _2273_ _2317_ _2319_ dmmu0.page_table\[14\]\[5\] _2325_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5051__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6723_ _0296_ clknet_leaf_44_core_clock dmmu0.page_table\[3\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3062__A1 net228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3935_ _1502_ _1596_ _1598_ _1599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_30_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinterconnect_inner_706 c0_i_core_int_sreg[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_34_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinterconnect_inner_717 c0_i_core_int_sreg[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_74_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinterconnect_inner_728 c1_i_core_int_sreg[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_74_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6654_ _0227_ clknet_leaf_31_core_clock dmmu0.page_table\[11\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3866_ _1525_ _1527_ _1529_ _1531_ _1532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_46_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5605_ _2690_ _0324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_41_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6585_ _0158_ clknet_leaf_18_core_clock immu_0.page_table\[3\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3797_ _1391_ _1462_ _1464_ _1465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input186_I c1_sr_bus_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3996__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3365__A2 _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5536_ _2651_ _0294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_83_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6572__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5467_ immu_1.high_addr_off\[7\] _1864_ _2603_ _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3165__I net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput630 net630 ic1_mem_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_30_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput641 net641 ic1_wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_44_1058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input353_I ic1_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput652 net652 ic1_wb_i_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5511__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4418_ _1769_ _1788_ _1975_ _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_4
Xoutput663 net663 inner_wb_adr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_61_2084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput674 net674 inner_wb_adr[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5398_ _1785_ _2570_ _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_1481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input47_I c0_o_mem_high_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput685 net685 inner_wb_o_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput696 net696 inner_wb_o_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7137_ net75 net599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4349_ _1858_ _1927_ _1929_ net1008 _1935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_35_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6067__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7068_ net407 net465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4617__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5814__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6019_ _2786_ _2924_ _2926_ dmmu1.page_table\[3\]\[3\] _2930_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3053__A1 net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3784__B _1452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3276__S _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5750__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4305__A1 net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4856__A2 _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5656__I1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3816__B1 _1473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_2075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3292__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5408__I1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6445__CLK clknet_leaf_26_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5569__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5033__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_2015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_2026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5666__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ net313 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_71_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3595__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4792__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6595__CLK clknet_leaf_24_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3651_ _1329_ _1330_ _1331_ net671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_77_2534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4544__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _0752_ clknet_leaf_71_core_clock immu_1.page_table\[12\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_2409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3582_ _1291_ net424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_1481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5321_ _2463_ _2516_ _2518_ dmmu0.page_table\[12\]\[7\] _2526_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5252_ _2485_ _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_48_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4847__A2 _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4203_ _1769_ _1834_ _1837_ _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_4
XANTENNA__3713__I _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5183_ _2441_ _0151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6049__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4134_ net83 net76 _1780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_3_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4065_ _1712_ _1713_ _1718_ _1724_ _0813_ _1725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_39_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3283__A1 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input101_I c0_sr_bus_data_o[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6938__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4967_ _2314_ _0062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_43_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3130__S1 _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3918_ net7 immu_0.high_addr_off\[2\] _1581_ _1582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_6706_ _0279_ clknet_leaf_98_core_clock dmmu0.page_table\[4\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4898_ _1802_ _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_85_1114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6637_ _0210_ clknet_leaf_11_core_clock dmmu0.page_table\[12\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3849_ immu_1.page_table\[12\]\[4\] immu_1.page_table\[13\]\[4\] immu_1.page_table\[14\]\[4\]
+ immu_1.page_table\[15\]\[4\] _1441_ _1442_ _1515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3096__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5732__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6568_ _0141_ clknet_leaf_21_core_clock immu_0.page_table\[5\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5519_ _2527_ _2630_ _2632_ net1077 _2641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6499_ _0072_ clknet_leaf_28_core_clock dmmu0.page_table\[14\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_37_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4299__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput460 net460 c0_i_req_data_valid vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput471 net471 c1_i_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput482 net482 c1_i_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput493 net493 c1_i_req_data[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6468__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_28_core_clock_I clknet_4_5__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5263__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3274__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4471__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5015__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3577__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5971__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4829__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3188__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_85_2803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3689__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3265__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5870_ _2790_ _2836_ _2838_ net886 _2844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4821_ _2221_ _0009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4752_ _2181_ _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4765__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3703_ immu_0.page_table\[12\]\[0\] immu_0.page_table\[13\]\[0\] immu_0.page_table\[14\]\[0\]
+ immu_0.page_table\[15\]\[0\] _1370_ _1372_ _1373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA_clkbuf_leaf_30_core_clock_I clknet_4_5__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4683_ _1839_ _2137_ _2138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3708__I _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6422_ _0804_ clknet_leaf_111_core_clock immu_0.page_table\[12\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4517__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3634_ _1320_ net687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4517__B2 dmmu1.page_table\[14\]\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5714__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5190__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6353_ _0735_ clknet_leaf_78_core_clock immu_1.page_table\[13\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3565_ net212 _1204_ _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_64_1754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5304_ _2515_ _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_64_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6284_ _0666_ clknet_leaf_39_core_clock dmmu0.page_table\[0\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3496_ net51 dmmu0.long_off_reg\[6\] _1234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5235_ _2476_ _0168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6610__CLK clknet_leaf_17_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5493__A2 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input149_I c1_o_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5166_ _2258_ _2430_ _2432_ net749 _2433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4117_ _1764_ _1768_ _1771_ net684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5097_ _2275_ _2382_ _2384_ immu_0.page_table\[7\]\[6\] _2391_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input316_I ic0_wb_adr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4048_ net11 immu_0.high_addr_off\[6\] _1708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3256__A1 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_26_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5999_ _2847_ _2907_ _2909_ dmmu1.page_table\[4\]\[8\] _2918_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_23_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5953__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3554__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3781__C _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6290__CLK clknet_leaf_101_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3495__A1 net51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4692__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold9 dmmu0.page_table\[2\]\[1\] net743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5236__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3247__A1 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3098__I1 net26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3342__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_46_core_clock clknet_4_13__leaf_core_clock clknet_leaf_46_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_70_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4747__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3528__I _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3972__B net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5172__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6633__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_96_core_clock_I clknet_4_9__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3350_ _0894_ _1083_ _1092_ _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_1938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6121__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3281_ dmmu0.page_table\[10\]\[4\] dmmu0.page_table\[11\]\[4\] _0865_ _1027_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5475__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5020_ _2346_ _0083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_85_core_clock clknet_4_10__leaf_core_clock clknet_leaf_85_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3089__I1 net22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6971_ _0544_ clknet_leaf_62_core_clock dmmu1.page_table\[0\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4435__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5922_ _2874_ _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4986__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5853_ _2833_ _0429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4804_ _1800_ _2208_ _2210_ immu_0.page_table\[13\]\[2\] _2213_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5935__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5784_ _2794_ _2778_ _2780_ net757 _2795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4202__A3 _1836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4735_ _2169_ _0784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3410__A1 _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ _2061_ _2123_ _2125_ net939 _2129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6405_ _0787_ clknet_leaf_1_core_clock immu_0.page_table\[14\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3617_ _1308_ net265 _1312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_4_9__f_core_clock clknet_3_4_0_core_clock clknet_4_9__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4597_ _1868_ _2075_ _2077_ net993 _2087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_40_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input266_I dcache_wb_o_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6336_ _0718_ clknet_leaf_78_core_clock immu_1.page_table\[15\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3548_ net136 net31 _1267_ _1274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6267_ _0649_ clknet_leaf_89_core_clock immu_1.page_table\[4\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3479_ _1209_ _1214_ _1217_ _1051_ _1218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5218_ _2465_ _0162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6198_ _0580_ clknet_leaf_5_core_clock immu_0.page_table\[11\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4674__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5149_ _2273_ _2414_ _2416_ net1092 _2422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3324__S1 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6506__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4044__I3 _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output485_I net485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6656__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4179__I net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6103__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4907__I _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5209__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4968__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_1562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4520_ _2039_ _0699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold206 dmmu0.page_table\[2\]\[7\] net940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4451_ _1996_ _1978_ _1981_ dmmu0.page_table\[0\]\[12\] _1997_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5145__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold217 dmmu1.page_table\[4\]\[9\] net951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold228 immu_1.page_table\[10\]\[7\] net962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3402_ net49 dmmu0.long_off_reg\[4\] _1142_ _1143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5696__A2 _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold239 dmmu1.page_table\[2\]\[11\] net973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7170_ net169 net625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4382_ _1953_ _0647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3207__B _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6121_ _2849_ _2975_ _2977_ dmmu1.page_table\[0\]\[9\] _2987_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3333_ net45 dmmu0.long_off_reg\[0\] _1077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_42_1145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6052_ _2948_ _0513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_7_Right_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3459__A1 _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3264_ _0889_ _1008_ _1009_ _0931_ _1010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_5003_ _1790_ _2222_ _2336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4120__A2 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3721__I _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3195_ dmmu0.page_table\[0\]\[1\] dmmu0.page_table\[1\]\[1\] dmmu0.page_table\[2\]\[1\]
+ dmmu0.page_table\[3\]\[1\] _0864_ _0867_ _0944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6529__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6954_ _0527_ clknet_leaf_57_core_clock dmmu1.page_table\[1\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5905_ _2792_ _2856_ _2858_ dmmu1.page_table\[7\]\[6\] _2865_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3631__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6885_ _0458_ clknet_leaf_55_core_clock dmmu1.page_table\[6\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6679__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5836_ _1802_ _2819_ _2821_ net1009 _2825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_57_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5384__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5767_ _2783_ _0393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input383_I ic1_wb_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4718_ _1797_ _2157_ _2159_ immu_0.page_table\[15\]\[1\] _2161_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5698_ _1892_ _2028_ _2031_ _2742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA_input77_I c0_sr_bus_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4649_ _2118_ _0749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_2066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6319_ _0701_ clknet_leaf_71_core_clock dmmu1.page_table\[14\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4111__A2 net379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7103__I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_2020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3870__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3481__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_1877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3806__I _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5678__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3233__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3689__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4102__A2 net326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3541__I _1270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput360 ic1_mem_data[7] net360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput371 ic1_wb_adr[2] net371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput382 ic1_wb_stb net382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_19_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5850__A2 _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput393 inner_wb_i_dat[13] net393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3861__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6821__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5063__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5602__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3951_ net112 immu_1.high_addr_off\[2\] _1614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3613__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4810__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6670_ _0243_ clknet_leaf_103_core_clock immu_0.high_addr_off\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3882_ net110 immu_1.high_addr_off\[0\] _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5621_ _2698_ _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4169__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6971__CLK clknet_leaf_62_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5552_ _2659_ _0302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4503_ _1870_ _2013_ _2015_ immu_1.page_table\[3\]\[10\] _2027_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5118__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5483_ _2459_ _2613_ _2615_ net968 _2621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6201__CLK clknet_leaf_103_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4434_ _1987_ _0665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3224__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7153_ net393 net608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4341__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4365_ _1824_ _1942_ _1944_ net963 _1945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_1674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6104_ _2978_ _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3316_ _1054_ _1056_ _1058_ _1060_ _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_61_1598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7084_ net337 net490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_67_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4296_ _1903_ _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6035_ net199 _2923_ _2925_ dmmu1.page_table\[3\]\[11\] _2938_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_52_1772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3247_ _0889_ _0991_ _0992_ _0902_ _0993_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_52_1783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input131_I c1_o_mem_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input229_I dcache_mem_o_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3178_ dmmu1.page_table\[0\]\[1\] dmmu1.page_table\[1\]\[1\] dmmu1.page_table\[2\]\[1\]
+ dmmu1.page_table\[3\]\[1\] _0888_ _0910_ _0927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_55_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6937_ _0510_ clknet_leaf_56_core_clock dmmu1.page_table\[2\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4282__I _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6868_ _0441_ clknet_leaf_67_core_clock dmmu1.page_table\[8\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_46_1587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_2081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5819_ _2814_ _0414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6799_ _0372_ clknet_leaf_66_core_clock dmmu1.page_table\[12\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3215__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4868__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output448_I net448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6085__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3518__S1 net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4096__A1 _1747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6844__CLK clknet_leaf_68_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5293__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3843__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5045__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5596__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4399__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6994__CLK clknet_leaf_97_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5348__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5899__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4020__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3454__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_35_core_clock_I clknet_4_7__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4571__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6374__CLK clknet_leaf_73_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_2337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4323__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_2348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4150_ _1795_ _0573_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3101_ _0853_ net540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4081_ _1502_ _1735_ _1740_ _1408_ _1741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4087__A1 net12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3032_ inner_wb_arbiter.o_sel_sig _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_37_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput190 c1_sr_bus_addr[3] net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_69_2277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5587__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4983_ _2324_ _0068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_2065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6722_ _0295_ clknet_leaf_39_core_clock dmmu0.page_table\[3\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3934_ _1434_ _1597_ _1598_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3062__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinterconnect_inner_707 c0_i_core_int_sreg[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_inner_718 c0_i_core_int_sreg[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_inner_729 c1_i_core_int_sreg[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_15_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3865_ _1375_ _1530_ _1383_ _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6653_ _0226_ clknet_leaf_17_core_clock dmmu0.page_table\[11\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5604_ _2459_ _2681_ _2684_ net930 _2690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_41_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3796_ _1463_ immu_0.page_table\[15\]\[2\] _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_41_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6584_ _0157_ clknet_leaf_24_core_clock immu_0.page_table\[3\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6717__CLK clknet_leaf_11_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5535_ _2451_ _2647_ _2649_ net1097 _2651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3996__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5466_ _2610_ _0265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input179_I c1_o_req_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput620 net620 ic1_mem_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput631 net631 ic1_mem_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput642 net642 ic1_wb_i_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_58_1970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4417_ _1974_ net91 _1784_ _1975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5511__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput653 net653 ic1_wb_i_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5397_ _1895_ net105 _2569_ _2570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput664 net664 inner_wb_adr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput675 net675 inner_wb_adr[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6867__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput686 net686 inner_wb_o_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input346_I ic1_mem_data[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput697 net697 inner_wb_o_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4348_ _1934_ _0632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7136_ net4 net598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4277__I _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6067__A2 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7067_ net407 net464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4279_ net188 net181 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
X_6018_ _2929_ _0498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_1810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5814__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6247__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3053__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4002__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6397__CLK clknet_leaf_112_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3436__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output565_I net565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5750__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3816__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5569__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_2005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_2027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3650_ _1306_ net242 _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_2524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3581_ net227 _1204_ _1291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_49_1460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5320_ _2525_ _0204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5251_ _1789_ _2484_ _2485_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_80_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4202_ net210 _1835_ _1836_ _1837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5182_ _2328_ _2430_ _2432_ net901 _2441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6049__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4133_ _1778_ net84 _1779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_3_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5257__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4064_ _1382_ _1723_ _1724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_30_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4966_ _1994_ _2298_ _2301_ dmmu0.page_table\[7\]\[11\] _2314_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6705_ _0278_ clknet_leaf_70_core_clock dmmu0.page_table\[4\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3917_ _1553_ _1554_ _1580_ _1581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_7_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4897_ _2268_ _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4560__I _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input296_I ic0_mem_data[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6636_ _0209_ clknet_leaf_13_core_clock dmmu0.page_table\[12\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3848_ _1514_ net666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5732__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3779_ immu_1.page_table\[12\]\[1\] immu_1.page_table\[13\]\[1\] immu_1.page_table\[14\]\[1\]
+ immu_1.page_table\[15\]\[1\] _1441_ _1442_ _1448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_6567_ _0140_ clknet_leaf_26_core_clock immu_0.page_table\[5\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5518_ _2640_ _0287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_56_1907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6498_ _0071_ clknet_leaf_32_core_clock dmmu0.page_table\[14\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_37_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput450 net450 c0_i_req_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5449_ net191 _1836_ _2600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4299__A1 _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput461 net461 c0_rst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_30_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput472 net472 c1_i_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput483 net483 c1_i_mem_exception vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput494 net494 c1_i_req_data[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_61_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7119_ net395 net572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_3_5_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7111__I net402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4471__A1 _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_36_core_clock clknet_4_7__leaf_core_clock clknet_leaf_36_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5420__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output682_I net682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4774__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5971__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3409__S0 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3086__I _0845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5487__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6412__CLK clknet_leaf_112_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3352__I3 dmmu0.page_table\[7\]\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_75_core_clock clknet_4_11__leaf_core_clock clknet_leaf_75_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_85_2804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6562__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4820_ _1821_ _2207_ _2209_ net1019 _2221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4751_ _1803_ _2175_ _2177_ immu_0.page_table\[14\]\[3\] _2181_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4765__A2 _2174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3702_ _1371_ _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_12_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4682_ _1826_ _1909_ _2137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_50_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3633_ _0812_ net258 _1320_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6421_ _0803_ clknet_leaf_1_core_clock immu_0.page_table\[12\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4517__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5714__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4073__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3564_ _1218_ _1281_ _1282_ net533 net542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6352_ _0734_ clknet_leaf_72_core_clock immu_1.page_table\[13\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5303_ _1977_ _2189_ _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6283_ _0665_ clknet_leaf_39_core_clock dmmu0.page_table\[0\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3495_ net51 dmmu0.long_off_reg\[6\] _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6100__I _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5234_ _2455_ _2470_ _2472_ immu_0.page_table\[2\]\[3\] _2476_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_1452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5165_ _2431_ _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4116_ _1770_ _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_58_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ _2390_ _0115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4047_ _1306_ _1696_ _1706_ _1707_ net673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_49_1700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__A1 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input211_I core_reset vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input309_I ic0_wb_adr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4205__A1 _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5998_ _2917_ _0490_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5953__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4949_ _2305_ _0053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_1855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6619_ _0192_ clknet_leaf_24_core_clock immu_0.page_table\[0\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_1699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6435__CLK clknet_leaf_112_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7106__I net397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6010__I _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6130__A1 net559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_58_Left_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output528_I net528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4692__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3878__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_2057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_4__f_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Left_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4747__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3558__I0 net160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5172__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3802__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_76_Left_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6121__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3280_ _0948_ _1022_ _1025_ _0875_ _1026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_29_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6928__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4683__A1 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5880__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6970_ _0543_ clknet_leaf_62_core_clock dmmu1.page_table\[0\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4435__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5921_ _1770_ _2872_ _2874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4986__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_85_Left_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5852_ net94 _2818_ _2820_ dmmu0.page_table\[1\]\[11\] _2833_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6308__CLK clknet_leaf_89_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4803_ _2212_ _0000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5935__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5783_ _1863_ _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_84_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4734_ _1819_ _2157_ _2159_ immu_0.page_table\[15\]\[9\] _2169_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4665_ _2128_ _0755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6458__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6404_ _0786_ clknet_leaf_110_core_clock immu_0.page_table\[14\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3616_ _1311_ net693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4596_ _2086_ _0728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4371__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6335_ _0717_ clknet_leaf_77_core_clock immu_1.page_table\[15\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3547_ _1273_ net544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input161_I c1_o_mem_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input259_I dcache_wb_o_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6266_ _0648_ clknet_leaf_86_core_clock immu_1.page_table\[4\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3478_ net156 dmmu1.long_off_reg\[6\] _1216_ _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5217_ _2328_ _2447_ _2449_ immu_0.page_table\[3\]\[8\] _2465_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4674__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6197_ _0579_ clknet_leaf_6_core_clock immu_0.page_table\[11\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5148_ _2421_ _0136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input22_I c0_o_mem_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5079_ _2332_ _2366_ _2368_ immu_0.page_table\[8\]\[10\] _2380_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output478_I net478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6103__A1 _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5862__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3313__B _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4968__A2 _2298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5917__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3539__I _1269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6600__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4028__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4450_ net95 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5145__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold207 dmmu1.page_table\[8\]\[0\] net941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold218 dmmu0.page_table\[3\]\[3\] net952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6750__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold229 immu_1.page_table\[4\]\[0\] net963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3401_ _1140_ _1122_ _1141_ _1142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4353__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4381_ _1866_ _1942_ _1944_ net877 _1953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3332_ _1072_ _1073_ _1074_ _1075_ _0877_ _0878_ _1076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_6120_ _2986_ _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6051_ _2788_ _2941_ _2943_ dmmu1.page_table\[2\]\[4\] _2948_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3263_ _0899_ dmmu1.page_table\[12\]\[4\] _1009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_1591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4656__A1 _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5002_ _2335_ _0076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3194_ _0940_ _0942_ _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4120__A3 _0815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_42_core_clock_I clknet_4_12__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6953_ _0526_ clknet_leaf_58_core_clock dmmu1.page_table\[1\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5904_ _2864_ _0449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6884_ _0457_ clknet_leaf_51_core_clock dmmu1.page_table\[6\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3631__A2 net257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5835_ _2824_ _0420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6280__CLK clknet_leaf_40_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5766_ _2782_ _2778_ _2780_ net868 _2783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5384__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3395__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4717_ _2160_ _0775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5697_ _2741_ _0365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input376_I ic1_wb_adr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4648_ _2069_ _2108_ _2110_ net982 _2118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4579_ _2051_ _2075_ _2077_ immu_1.page_table\[14\]\[0\] _2078_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6318_ _0700_ clknet_leaf_71_core_clock dmmu1.page_table\[14\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6249_ _0631_ clknet_leaf_90_core_clock immu_1.page_table\[5\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5844__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3870__A2 net238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6623__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output595_I net595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6021__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3386__A1 net153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4583__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3481__S1 _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6175__I1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3094__I _0849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3233__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3689__A2 net310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_1780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4638__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput350 ic1_mem_data[27] net350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput361 ic1_mem_data[8] net361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput372 ic1_wb_adr[3] net372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_1805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput383 ic1_wb_we net383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput394 inner_wb_i_dat[14] net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_19_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold90 dmmu0.page_table\[1\]\[2\] net824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3861__A2 _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5063__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_2050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3950_ net112 immu_1.high_addr_off\[2\] _1613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3613__A2 net263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4810__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3881_ _1502_ _1539_ _1545_ _1408_ _1546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_2_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5620_ _1976_ _2412_ _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_39_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3377__A1 net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5551_ _2529_ _2647_ _2649_ net772 _2659_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4502_ _2026_ _0694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5118__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5482_ _2620_ _0271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3218__B _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4433_ _1806_ _1979_ _1982_ dmmu0.page_table\[0\]\[4\] _1987_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3224__S1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7152_ net392 net607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4364_ _1943_ _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6079__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6103_ _1823_ _2975_ _2977_ net981 _2978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3315_ _0938_ _1059_ _1060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7083_ net336 net489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4295_ _1857_ _1894_ _1897_ immu_1.page_table\[0\]\[5\] _1903_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6034_ _2937_ _0506_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3246_ _0908_ dmmu1.page_table\[4\]\[4\] _0992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_52_1773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3301__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3177_ _0897_ _0925_ _0926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6646__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input124_I c1_o_mem_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4563__I _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6936_ _0509_ clknet_leaf_56_core_clock dmmu1.page_table\[2\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6867_ _0440_ clknet_leaf_45_core_clock dmmu1.page_table\[8\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5818_ _2103_ _2802_ _2804_ net816 _2814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6798_ _0371_ clknet_leaf_53_core_clock dmmu1.page_table\[12\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_1108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5749_ _2771_ _0387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4317__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3215__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4868__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4738__I net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7114__I net390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5293__A1 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output510_I net510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5045__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5596__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_2080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5348__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3359__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3454__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_2463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6669__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5808__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3100_ net132 net27 _0850_ _0853_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4080_ _1502_ _1737_ _1739_ _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_37_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3031_ _0811_ net559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_56_1602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput180 c1_o_req_ppl_submit net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput191 c1_sr_bus_addr[4] net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_69_2278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3390__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4982_ _2271_ _2317_ _2319_ dmmu0.page_table\[14\]\[4\] _2324_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5587__A2 _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6721_ _0294_ clknet_leaf_41_core_clock dmmu0.page_table\[3\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3933_ immu_1.page_table\[12\]\[6\] immu_1.page_table\[13\]\[6\] immu_1.page_table\[14\]\[6\]
+ immu_1.page_table\[15\]\[6\] _1474_ _1433_ _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_50_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_inner_708 c0_i_core_int_sreg[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_6652_ _0225_ clknet_leaf_28_core_clock dmmu0.page_table\[11\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinterconnect_inner_719 c0_i_core_int_sreg[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_3864_ immu_0.page_table\[12\]\[4\] immu_0.page_table\[13\]\[4\] immu_0.page_table\[14\]\[4\]
+ immu_0.page_table\[15\]\[4\] _1463_ _1371_ _1530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_73_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5603_ _2689_ _0323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6583_ _0156_ clknet_leaf_24_core_clock immu_0.page_table\[3\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_41_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3795_ _1369_ _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_6_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6199__CLK clknet_leaf_6_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5534_ _2650_ _0293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5465_ immu_1.high_addr_off\[6\] _1861_ _2603_ _2610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput610 net610 ic0_wb_i_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_23_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput621 net621 ic1_mem_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput632 net632 ic1_mem_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4416_ net90 _1974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
Xoutput643 net643 ic1_wb_i_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5511__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput654 net654 ic1_wb_i_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput665 net665 inner_wb_adr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5396_ net86 _1787_ _1971_ _1972_ _2569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_41_1915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput676 net676 inner_wb_adr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3522__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput687 net687 inner_wb_o_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7135_ net65 net588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4347_ _1855_ _1927_ _1929_ immu_1.page_table\[5\]\[4\] _1934_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput698 net698 inner_wb_o_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input241_I dcache_wb_adr[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Left_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_35_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input339_I ic1_mem_data[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7066_ net406 net463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4278_ _1872_ _1825_ _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__5275__A1 net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6017_ _2784_ _2924_ _2926_ net928 _2929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3229_ dmmu0.page_table\[0\]\[3\] dmmu0.page_table\[1\]\[3\] dmmu0.page_table\[2\]\[3\]
+ dmmu0.page_table\[3\]\[3\] _0950_ _0952_ _0976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_39_1866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5027__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3411__B _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_26_core_clock clknet_4_5__leaf_core_clock clknet_leaf_26_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_1167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3589__A1 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4786__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6919_ _0492_ clknet_leaf_60_core_clock dmmu1.page_table\[4\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4250__A2 net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Left_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4002__A2 _1663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7109__I net400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3436__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5750__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3761__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6811__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_2104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_65_core_clock clknet_4_15__leaf_core_clock clknet_leaf_65_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6961__CLK clknet_leaf_64_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_2044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3816__A2 _1459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_2710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_2721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_2131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5569__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_2153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3124__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_2006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_2075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6341__CLK clknet_leaf_73_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4529__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3547__I _1273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_2514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_2042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_2525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3201__B1 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3580_ _1290_ net423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3991__B net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3752__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_1325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6491__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5250_ _1971_ _2205_ _2484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_23_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4201_ net194 net193 net192 _1836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_62_1683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5181_ _2440_ _0150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4132_ net85 _1778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_3_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5257__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4063_ _1378_ _1720_ _1722_ _1723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_30_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5009__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4965_ _2313_ _0061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_43_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6704_ _0277_ clknet_leaf_99_core_clock dmmu0.page_table\[4\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3916_ net6 immu_0.high_addr_off\[1\] _1580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4896_ _2267_ _2261_ _2263_ net933 _2268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6635_ _0208_ clknet_leaf_12_core_clock dmmu0.page_table\[12\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3847_ net237 _1513_ _1360_ _1514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6834__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input191_I c1_sr_bus_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input289_I ic0_mem_data[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6566_ _0139_ clknet_leaf_22_core_clock immu_0.page_table\[5\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5732__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3778_ _1440_ _1443_ _1444_ _1445_ _1446_ _1447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_6_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5517_ _2463_ _2630_ _2632_ dmmu0.page_table\[13\]\[7\] _2640_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_1425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6497_ _0070_ clknet_leaf_16_core_clock dmmu0.page_table\[14\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_37_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5448_ _1895_ net210 _2599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input52_I c0_o_mem_high_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput440 net440 c0_i_req_data[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4299__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput451 net451 c0_i_req_data[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput462 net462 c1_disable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6984__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput473 net473 c1_i_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput484 net484 c1_i_req_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3192__I _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5379_ _2560_ _0228_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput495 net495 c1_i_req_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7118_ net394 net571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5248__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6214__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7049_ net285 net436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_29_Right_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3354__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_2108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4471__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6364__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4759__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5420__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5971__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3982__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Right_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3409__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5184__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4931__B1 _2291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_2081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5487__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_47_Right_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_66_2204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6707__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_47_core_clock_I clknet_4_13__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6857__CLK clknet_leaf_101_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4750_ _2180_ _0788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_1936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_56_Right_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3701_ net313 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_3_1160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4681_ _2136_ _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6420_ _0802_ clknet_leaf_0_core_clock immu_0.page_table\[12\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3632_ _1319_ net686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5714__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4073__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3725__A1 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6351_ _0733_ clknet_leaf_72_core_clock immu_1.page_table\[13\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3563_ _1154_ _1186_ _1231_ _1282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_84_1171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5302_ _2514_ _0197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6282_ _0664_ clknet_leaf_40_core_clock dmmu0.page_table\[0\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3494_ _1204_ _1218_ _1232_ net532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_80_1068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6237__CLK clknet_leaf_95_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5233_ _2475_ _0167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_65_Right_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5164_ _1980_ _2429_ _2431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4115_ _1769_ _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5095_ _2273_ _2382_ _2384_ immu_0.page_table\[7\]\[5\] _2390_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6387__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4046_ _1535_ net244 _1707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4453__A2 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input204_I c1_sr_bus_data_o[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_74_Right_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4205__A2 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5997_ _2794_ _2907_ _2909_ dmmu1.page_table\[4\]\[7\] _2917_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_1560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4948_ _2267_ _2299_ _2302_ net740 _2305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5953__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3964__A1 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4879_ _2255_ _0033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_1867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5166__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6618_ _0191_ clknet_leaf_19_core_clock immu_0.page_table\[0\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4913__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6549_ _0122_ clknet_leaf_9_core_clock immu_0.page_table\[6\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3915__I net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Right_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5469__A1 _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3851__S _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4692__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7122__I net67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3878__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_112_core_clock clknet_4_0__leaf_core_clock clknet_leaf_112_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1092 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3097__I _0851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5157__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3558__I1 net55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3802__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6121__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4683__A2 _2137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5880__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7032__I net277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__A1 _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4435__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5920_ _2872_ _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_0_13 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_3_0_core_clock clknet_0_core_clock clknet_3_3_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_17_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5851_ _2832_ _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4802_ _1797_ _2208_ _2210_ immu_0.page_table\[13\]\[1\] _2212_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5782_ _2793_ _0398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5935__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3946__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4733_ _2168_ _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4664_ _2059_ _2123_ _2125_ net761 _2128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6403_ _0785_ clknet_leaf_108_core_clock immu_0.page_table\[15\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3615_ _1308_ net264 _1311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3735__I _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4595_ _1866_ _2075_ _2077_ net810 _2086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_2107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4371__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6334_ _0716_ clknet_leaf_77_core_clock immu_1.page_table\[15\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3546_ net135 net30 _1267_ _1273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6265_ _0647_ clknet_leaf_87_core_clock immu_1.page_table\[4\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3477_ _1187_ _1190_ _1215_ _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5950__I _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input154_I c1_o_mem_high_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5216_ _2464_ _0161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6196_ _0578_ clknet_leaf_0_core_clock immu_0.page_table\[11\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4674__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4566__I _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5147_ _2271_ _2414_ _2416_ net764 _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_2058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input321_I ic0_wb_adr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5078_ _2379_ _0108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input15_I c0_o_mem_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4029_ _1439_ _1689_ _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3937__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6402__CLK clknet_leaf_112_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5139__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7117__I net393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6103__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5311__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5614__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5465__I1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5378__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3928__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4028__S1 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3555__I _1277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold208 immu_1.page_table\[8\]\[3\] net942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold219 dmmu0.page_table\[11\]\[2\] net953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3400_ net48 dmmu0.long_off_reg\[3\] _1141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4353__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4380_ _1952_ _0646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_1715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3331_ dmmu0.page_table\[8\]\[6\] dmmu0.page_table\[9\]\[6\] dmmu0.page_table\[10\]\[6\]
+ dmmu0.page_table\[11\]\[6\] _0864_ _0941_ _1075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_26_1879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4105__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6050_ _2947_ _0512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3262_ dmmu1.page_table\[13\]\[4\] _1008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input7_I c0_o_instr_long_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ _1996_ _2316_ _2318_ net1071 _2335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4656__A2 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3193_ dmmu0.page_table\[4\]\[1\] dmmu0.page_table\[5\]\[1\] dmmu0.page_table\[6\]\[1\]
+ dmmu0.page_table\[7\]\[1\] _0864_ _0941_ _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_56_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6952_ _0525_ clknet_leaf_54_core_clock dmmu1.page_table\[1\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5903_ _2790_ _2856_ _2858_ dmmu1.page_table\[7\]\[5\] _2864_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_2097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6883_ _0456_ clknet_leaf_68_core_clock dmmu1.page_table\[7\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6425__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5834_ _1799_ _2819_ _2821_ net824 _2824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5765_ _1845_ _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4716_ _1777_ _2157_ _2159_ immu_0.page_table\[15\]\[0\] _2160_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3395__A2 _1131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5696_ _2049_ _2725_ _2727_ dmmu1.page_table\[13\]\[12\] _2741_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6575__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4647_ _2117_ _0748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3465__I _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input271_I dcache_wb_o_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_1913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input369_I ic1_wb_adr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5541__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4578_ _2076_ _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6317_ _0699_ clknet_leaf_70_core_clock dmmu1.page_table\[14\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3529_ net142 net37 _0850_ _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_1247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6097__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6248_ _0630_ clknet_leaf_90_core_clock immu_1.page_table\[5\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5844__A1 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6179_ dmmu1.long_off_reg\[4\] _1855_ _3016_ _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_2077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6021__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output490_I net490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output588_I net588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4583__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4335__A1 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_1158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5590__I _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput340 ic1_mem_data[18] net340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3846__B1 _1503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput351 ic1_mem_data[28] net351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_1776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput362 ic1_mem_data[9] net362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput373 ic1_wb_adr[4] net373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold80 dmmu0.page_table\[13\]\[1\] net814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput384 inner_disable net384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput395 inner_wb_i_dat[15] net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xhold91 immu_1.page_table\[12\]\[0\] net825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_56_1828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6448__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5063__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3074__A1 net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4271__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4810__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3880_ _1502_ _1542_ _1544_ _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_85_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5765__I _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5550_ _2658_ _0301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4501_ _1868_ _2014_ _2016_ immu_1.page_table\[3\]\[9\] _2026_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5481_ _2457_ _2613_ _2615_ dmmu0.page_table\[4\]\[4\] _2620_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4432_ _1986_ _0664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5523__B1 _2631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7151_ net391 net606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4363_ _1912_ _1941_ _1943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6079__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6102_ _2976_ _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3314_ dmmu0.page_table\[4\]\[5\] dmmu0.page_table\[5\]\[5\] dmmu0.page_table\[6\]\[5\]
+ dmmu0.page_table\[7\]\[5\] _0872_ _0941_ _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_10_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7082_ net335 net488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4294_ _1902_ _0610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5826__A1 _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6033_ _2851_ _2923_ _2925_ net1104 _2937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3245_ dmmu1.page_table\[5\]\[4\] _0991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_52_1774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3176_ dmmu1.page_table\[4\]\[1\] dmmu1.page_table\[5\]\[1\] dmmu1.page_table\[6\]\[1\]
+ dmmu1.page_table\[7\]\[1\] _0908_ _0910_ _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_74_1917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_16_core_clock clknet_4_6__leaf_core_clock clknet_leaf_16_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input117_I c1_o_instr_long_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6935_ _0508_ clknet_leaf_64_core_clock dmmu1.page_table\[3\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6866_ _0439_ clknet_leaf_66_core_clock dmmu1.page_table\[8\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6003__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5817_ _2813_ _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6797_ _0370_ clknet_leaf_47_core_clock dmmu1.page_table\[12\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5748_ _2101_ _2760_ _2762_ net742 _2771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input82_I c0_sr_bus_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5679_ _2732_ _0356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4317__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4868__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_55_core_clock clknet_4_15__leaf_core_clock clknet_leaf_55_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_73_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5293__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output503_I net503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3798__C _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7130__I net60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5045__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6740__CLK clknet_leaf_44_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_2660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3359__A2 _1101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6890__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_94_core_clock clknet_4_8__leaf_core_clock clknet_leaf_94_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_49_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4308__A1 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5505__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_2464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_2339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5808__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6270__CLK clknet_leaf_90_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3030_ _0809_ _0810_ mem_dcache_arb.transfer_active _0811_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_1584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput170 c1_o_req_addr[15] net170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput181 c1_sr_bus_addr[0] net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_56_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput192 c1_sr_bus_addr[5] net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_69_2279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7040__I net307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3390__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_1423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3047__A1 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_104_core_clock_I clknet_4_2__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4981_ _2323_ _0067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3932_ _1440_ _1595_ _1596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6720_ _0293_ clknet_leaf_38_core_clock dmmu0.page_table\[3\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_1967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6651_ _0224_ clknet_leaf_30_core_clock dmmu0.page_table\[11\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_inner_709 c0_i_core_int_sreg[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_3863_ _1368_ _1528_ _1529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5602_ _2457_ _2681_ _2684_ dmmu0.page_table\[6\]\[4\] _2689_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5744__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6582_ _0155_ clknet_leaf_19_core_clock immu_0.page_table\[3\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3794_ _1385_ immu_0.page_table\[14\]\[2\] _1462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5533_ _2444_ _2647_ _2649_ net990 _2650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_1705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5464_ _2609_ _0264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput600 net600 ic0_mem_req vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_44_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput611 net611 ic0_wb_i_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput622 net622 ic1_mem_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4415_ _1971_ _1972_ _1973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xoutput633 net633 ic1_mem_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_2065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_54_core_clock_I clknet_4_15__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5395_ _2568_ _0236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput644 net644 ic1_wb_i_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6613__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput655 net655 ic1_wb_i_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput666 net666 inner_wb_adr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput677 net677 inner_wb_adr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7134_ net64 net587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput688 net688 inner_wb_o_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4346_ _1933_ _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_39_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput699 net699 inner_wb_o_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_61_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7065_ net211 net461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4277_ _1823_ _1890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_35_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input234_I dcache_wb_adr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6016_ _2928_ _0497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3228_ dmmu0.page_table\[4\]\[3\] dmmu0.page_table\[5\]\[3\] dmmu0.page_table\[6\]\[3\]
+ dmmu0.page_table\[7\]\[3\] _0950_ _0952_ _0975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_78_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6763__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4483__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3159_ _0900_ _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_input401_I inner_wb_i_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5027__A2 _2336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3038__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3589__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4786__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6918_ _0491_ clknet_leaf_61_core_clock dmmu1.page_table\[4\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5983__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6849_ _0422_ clknet_leaf_37_core_clock dmmu0.page_table\[1\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwire705 _1407_ net705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_52_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3854__S _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output453_I net453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6293__CLK clknet_leaf_82_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7125__I net70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4710__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_5_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3816__A3 _1468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_2700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_2711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_1907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_2722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3124__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_2007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_60_2018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_2029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4529__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3201__A1 _0930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3201__B2 _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6636__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6151__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7035__I net302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4200_ net191 _1835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5180_ _2277_ _2430_ _2432_ immu_0.page_table\[4\]\[7\] _2440_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6786__CLK clknet_leaf_46_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4131_ _1776_ _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_3_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_2082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5257__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4062_ _1366_ _1721_ _1722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_30_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4465__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5009__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4217__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5965__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4964_ _1821_ _2298_ _2301_ dmmu0.page_table\[7\]\[10\] _2313_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_28_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6703_ _0276_ clknet_leaf_41_core_clock dmmu0.page_table\[4\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3915_ net2 _1579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_28_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4895_ _1799_ _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3440__A1 net50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3846_ _1422_ _1490_ _1498_ _1503_ _1512_ _1513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6634_ _0207_ clknet_leaf_14_core_clock dmmu0.page_table\[12\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_1128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3777_ _1415_ _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
X_6565_ _0138_ clknet_leaf_22_core_clock immu_0.page_table\[5\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input184_I c1_sr_bus_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5516_ _2639_ _0286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6496_ _0069_ clknet_leaf_28_core_clock dmmu0.page_table\[14\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_56_1909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5447_ net325 _1766_ _2598_ _1771_ _0258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput430 net430 c0_i_req_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_37_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput441 net441 c0_i_req_data[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input351_I ic1_mem_data[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput452 net452 c0_i_req_data[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput463 net463 c1_i_core_int_sreg[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput474 net474 c1_i_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5378_ _2457_ _2553_ _2555_ dmmu0.page_table\[11\]\[4\] _2560_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput485 net485 c1_i_req_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input45_I c0_o_mem_high_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput496 net496 c1_i_req_data[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_leaf_6_core_clock clknet_4_1__leaf_core_clock clknet_leaf_6_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7117_ net393 net570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4329_ _1866_ _1911_ _1914_ net776 _1923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5248__A2 _2469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7048_ net284 net435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_22_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3354__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4759__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_102_core_clock clknet_4_3__leaf_core_clock clknet_leaf_102_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5420__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_26_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6659__CLK clknet_leaf_26_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5708__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3982__A2 _1639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5184__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4931__A1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4931__B2 _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5487__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3498__A1 net52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_2009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_1289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_2806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3670__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3700_ _1369_ _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_50_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4680_ _2105_ _2122_ _2124_ immu_1.page_table\[11\]\[10\] _2136_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _0812_ net257 _1319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_10_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6350_ _0732_ clknet_leaf_63_core_clock immu_1.page_table\[13\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3562_ _1169_ _1202_ _1281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_45_1112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5301_ net93 _2501_ _2503_ immu_0.page_table\[0\]\[10\] _2514_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_80_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6281_ _0663_ clknet_leaf_39_core_clock dmmu0.page_table\[0\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3493_ _1219_ _1231_ _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5232_ _2453_ _2470_ _2472_ immu_0.page_table\[2\]\[2\] _2475_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3489__A1 net50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5163_ _2429_ _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4114_ net211 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5094_ _2389_ _0114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_1517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4045_ net2 _1700_ _1705_ _1382_ _1422_ _1706_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_49_1702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4453__A3 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3661__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6801__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5996_ _2916_ _0489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_26_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4947_ _2304_ _0052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input399_I inner_wb_i_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3964__A2 _1626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4878_ _1821_ _2241_ _2243_ dmmu0.page_table\[9\]\[10\] _2255_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6951__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5166__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6617_ _0190_ clknet_leaf_24_core_clock immu_0.page_table\[0\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3829_ _1372_ _1492_ _1495_ _1366_ _1496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_43_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4913__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6548_ _0121_ clknet_leaf_5_core_clock immu_0.page_table\[6\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6115__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6479_ _0052_ clknet_leaf_35_core_clock dmmu0.page_table\[7\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6331__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4429__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3652__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6481__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5929__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_2046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5157__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_3_1_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4668__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5880__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6824__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5093__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5768__I _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3643__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5850_ _2531_ _2818_ _2820_ net964 _2832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4801_ _2211_ _0808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5396__A1 net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6974__CLK clknet_leaf_64_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5781_ _2792_ _2778_ _2780_ net854 _2793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_1723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4732_ _1817_ _2157_ _2159_ immu_0.page_table\[15\]\[8\] _2168_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3946__A2 _1605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4663_ _2127_ _0754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6204__CLK clknet_leaf_97_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ _0784_ clknet_leaf_112_core_clock immu_0.page_table\[15\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3614_ _1310_ net692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4594_ _2085_ _0727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3237__B _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3545_ _1272_ net558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4371__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6333_ _0715_ clknet_leaf_76_core_clock immu_1.page_table\[15\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ _0646_ clknet_leaf_86_core_clock immu_1.page_table\[4\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3476_ net155 dmmu1.long_off_reg\[5\] _1215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6354__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5215_ _2463_ _2447_ _2449_ net1099 _2464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6195_ _0577_ clknet_leaf_4_core_clock immu_0.page_table\[11\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input147_I c1_o_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5146_ _2420_ _0135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5077_ _2330_ _2367_ _2369_ net980 _2379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input314_I ic0_wb_adr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4028_ immu_1.page_table\[8\]\[9\] immu_1.page_table\[9\]\[9\] immu_1.page_table\[10\]\[9\]
+ immu_1.page_table\[11\]\[9\] _1409_ _1410_ _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_79_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4831__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5979_ _1873_ _1892_ _2030_ _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_75_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5139__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output533_I net533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5311__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7133__I net63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6847__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5075__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5614__A2 _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3625__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6997__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3102__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_109_core_clock_I clknet_4_0__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5378__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6227__CLK clknet_leaf_90_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4050__A1 net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6377__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold209 dmmu0.page_table\[8\]\[7\] net943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4353__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3330_ dmmu0.page_table\[12\]\[6\] dmmu0.page_table\[13\]\[6\] dmmu0.page_table\[14\]\[6\]
+ dmmu0.page_table\[15\]\[6\] _0864_ _0941_ _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_21_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4105__A2 net381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3261_ _0889_ _1005_ _1006_ _1007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7043__I net279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_59_core_clock_I clknet_4_15__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5000_ _2334_ _0075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4656__A3 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3192_ _0867_ _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_59_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6951_ _0524_ clknet_leaf_53_core_clock dmmu1.page_table\[1\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5902_ _2863_ _0448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6882_ _0455_ clknet_leaf_66_core_clock dmmu1.page_table\[7\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5833_ _2823_ _0419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5764_ _2781_ _0392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4715_ _2158_ _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5695_ _2740_ _0364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4646_ _2067_ _2108_ _2110_ net1063 _2117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_12_Left_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5541__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4577_ _1912_ _2074_ _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_2085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input264_I dcache_wb_o_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_111_core_clock_I clknet_4_0__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6316_ _0698_ clknet_leaf_98_core_clock dmmu1.page_table\[14\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3528_ _1263_ net550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_45_core_clock clknet_4_12__leaf_core_clock clknet_leaf_45_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6097__A2 _2957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6247_ _0629_ clknet_leaf_87_core_clock immu_1.page_table\[5\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3459_ _0906_ _1198_ _1199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5844__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6178_ _3020_ _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _2409_ _0129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5402__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4804__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A1 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_61_core_clock_I clknet_4_14__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6021__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4032__A1 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3466__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4583__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7128__I net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_84_core_clock clknet_4_10__leaf_core_clock clknet_leaf_84_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4335__A2 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_1582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4099__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput330 ic1_mem_ack net330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3846__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput341 ic1_mem_data[19] net341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput352 ic1_mem_data[29] net352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput363 ic1_wb_adr[0] net363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput374 ic1_wb_adr[5] net374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold70 dmmu0.page_table\[8\]\[3\] net804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput385 inner_embed_mode net385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xhold81 dmmu1.page_table\[12\]\[8\] net815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput396 inner_wb_i_dat[1] net396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xhold92 dmmu1.page_table\[6\]\[8\] net826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_76_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3074__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4271__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7038__I net305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4500_ _2025_ _0693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5480_ _2619_ _0270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3209__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_1 _0847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4431_ _1803_ _1979_ _1982_ dmmu0.page_table\[0\]\[3\] _1986_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5523__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4362_ _1941_ _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7150_ net390 net605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6079__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6101_ _1770_ _2974_ _2976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3313_ _0940_ _1057_ _0958_ _1058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7081_ net334 net487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4293_ _1854_ _1894_ _1897_ immu_1.page_table\[0\]\[4\] _1902_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_43_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5287__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6032_ _2936_ _0505_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3244_ dmmu1.page_table\[6\]\[4\] dmmu1.page_table\[7\]\[4\] _0908_ _0990_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_52_1764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3175_ _0922_ _0923_ _0907_ _0924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5039__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6934_ _0507_ clknet_leaf_59_core_clock dmmu1.page_table\[3\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4065__C _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6542__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6865_ _0438_ clknet_leaf_46_core_clock dmmu1.page_table\[8\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6003__A2 _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5816_ _2101_ _2802_ _2804_ net1026 _2813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4014__A1 _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6796_ _0369_ clknet_leaf_48_core_clock dmmu1.page_table\[12\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1946 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5747_ _2770_ _0386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input381_I ic1_wb_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6692__CLK clknet_leaf_92_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5678_ _2061_ _2726_ _2728_ dmmu1.page_table\[13\]\[3\] _2732_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_33_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input75_I c0_o_req_ppl_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4317__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4629_ _2106_ _0741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3828__A1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4253__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_2650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4005__A1 net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6190__C _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_2093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_2590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5505__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4308__A2 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_2454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__CLK clknet_leaf_109_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5808__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput160 c1_o_mem_sel[0] net160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3295__A2 _1040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput171 c1_o_req_addr[1] net171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput182 c1_sr_bus_addr[10] net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput193 c1_sr_bus_addr[6] net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_1626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6565__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4980_ _2269_ _2317_ _2319_ net1087 _2323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3047__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3931_ immu_1.page_table\[8\]\[6\] immu_1.page_table\[9\]\[6\] immu_1.page_table\[10\]\[6\]
+ immu_1.page_table\[11\]\[6\] _1474_ _1433_ _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_74_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6650_ _0223_ clknet_leaf_10_core_clock dmmu0.page_table\[15\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3862_ immu_0.page_table\[8\]\[4\] immu_0.page_table\[9\]\[4\] immu_0.page_table\[10\]\[4\]
+ immu_0.page_table\[11\]\[4\] _1463_ _1391_ _1528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5601_ _2688_ _0322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5744__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6581_ _0154_ clknet_leaf_20_core_clock immu_0.page_table\[3\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3793_ immu_0.page_table\[12\]\[2\] immu_0.page_table\[13\]\[2\] _1396_ _1461_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5532_ _2648_ _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_42_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3850__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5463_ immu_1.high_addr_off\[5\] _1858_ _2603_ _2609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput601 net601 ic0_rst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_80_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput612 net612 ic0_wb_i_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4414_ net83 net76 _1972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xoutput623 net623 ic1_mem_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_58_1951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput634 net634 ic1_mem_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5394_ _1996_ _2552_ _2554_ net1074 _2568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput645 net645 ic1_wb_i_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput656 net656 ic1_wb_i_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_54_1826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7133_ net63 net586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput667 net667 inner_wb_adr[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4180__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput678 net678 inner_wb_adr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4345_ _1852_ _1927_ _1929_ immu_1.page_table\[5\]\[3\] _1933_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput689 net689 inner_wb_o_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7064_ net276 net460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4276_ _1889_ _0605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_35_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6908__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6015_ _2782_ _2924_ _2926_ net1051 _2928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3227_ _0883_ _0973_ _0879_ _0974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4855__I _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4483__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5680__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input227_I dcache_mem_o_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3158_ _0898_ _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_59_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3038__A2 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3089_ net127 net22 _0842_ _0847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5432__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6917_ _0490_ clknet_leaf_57_core_clock dmmu1.page_table\[4\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5983__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4786__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6848_ _0421_ clknet_leaf_48_core_clock dmmu0.page_table\[1\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6779_ _0352_ clknet_leaf_104_core_clock dmmu0.long_off_reg\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6438__CLK clknet_leaf_26_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold370 dmmu1.page_table\[3\]\[10\] net1104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_output446_I net446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4710__A2 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6588__CLK clknet_leaf_17_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7141__I net396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_2701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_2712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3029__A2 net159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_2144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_2008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_2019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_2090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4529__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5726__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_77_2516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_77_2538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3832__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6151__A1 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3780__S _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4130_ net92 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_20_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4061_ immu_0.page_table\[12\]\[10\] immu_0.page_table\[13\]\[10\] immu_0.page_table\[14\]\[10\]
+ immu_0.page_table\[15\]\[10\] _1487_ _1390_ _1721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_78_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4465__A1 _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7051__I net287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4217__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5965__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4963_ _2312_ _0060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_47_1641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6702_ _0275_ clknet_leaf_49_core_clock dmmu0.page_table\[4\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_28_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3914_ net659 _1577_ _1578_ net668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4894_ _2266_ _0037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6633_ _0206_ clknet_leaf_30_core_clock dmmu0.page_table\[12\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3845_ _0813_ _1511_ _1512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4076__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6564_ _0137_ clknet_leaf_27_core_clock immu_0.page_table\[5\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3776_ immu_1.page_table\[2\]\[1\] immu_1.page_table\[3\]\[1\] _1435_ _1445_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5515_ _2461_ _2630_ _2632_ net788 _2639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6495_ _0068_ clknet_leaf_32_core_clock dmmu0.page_table\[14\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input177_I c1_o_req_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5446_ _1422_ net379 _2598_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput420 net420 c0_i_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput431 net431 c0_i_req_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput442 net442 c0_i_req_data[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6730__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput453 net453 c0_i_req_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4153__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput464 net464 c1_i_core_int_sreg[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5377_ _2559_ _0227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput475 net475 c1_i_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input344_I ic1_mem_data[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput486 net486 c1_i_req_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7116_ net392 net569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput497 net497 c1_i_req_data[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_61_1184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4328_ _1922_ _0624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input38_I c0_o_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7047_ net283 net434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4259_ _1849_ _1876_ _1878_ immu_1.page_table\[7\]\[2\] _1881_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6880__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5410__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4759__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5708__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6260__CLK clknet_leaf_90_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5184__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output563_I net563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4931__A2 _2290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6040__I _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6133__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_0_Left_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_2807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3670__A2 net321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5947__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6603__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3630_ _1318_ net700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3186__A1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4383__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3561_ _1280_ net561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7046__I net282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5300_ _2513_ _0196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3507__C _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3492_ _0883_ _1223_ _1227_ _1230_ _1119_ _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_51_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6280_ _0662_ clknet_leaf_40_core_clock dmmu0.page_table\[0\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5231_ _2474_ _0166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4686__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5162_ _1789_ _2428_ _2429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4113_ net659 _1767_ _1768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5093_ _2271_ _2382_ _2384_ immu_0.page_table\[7\]\[4\] _2389_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4044_ _1701_ _1702_ _1703_ _1704_ _1367_ _1383_ _1705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__3110__A1 net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3661__A2 net373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5995_ _2792_ _2907_ _2909_ net920 _2916_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6283__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4946_ _2265_ _2299_ _2302_ dmmu0.page_table\[7\]\[1\] _2304_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_23_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3413__A2 _1153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_66_core_clock_I clknet_4_12__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4877_ _2254_ _0032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input294_I ic0_mem_data[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6616_ _0189_ clknet_leaf_17_core_clock immu_0.page_table\[0\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3828_ _1391_ _1493_ _1494_ _1495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5166__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3177__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6547_ _0120_ clknet_leaf_10_core_clock immu_0.page_table\[7\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4913__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3759_ immu_0.page_table\[6\]\[1\] immu_0.page_table\[7\]\[1\] immu_0.page_table\[14\]\[1\]
+ immu_0.page_table\[15\]\[1\] _1370_ _1377_ _1428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_28_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_18_Left_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6115__A1 _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6478_ _0051_ clknet_leaf_32_core_clock dmmu0.page_table\[7\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5429_ _2589_ _0249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_7_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5874__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4429__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5626__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_27_Left_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6626__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3652__A2 net371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5929__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_6__f_core_clock clknet_3_3_0_core_clock clknet_4_6__leaf_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_1769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4601__A1 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output680_I net680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6776__CLK clknet_leaf_104_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5157__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_36_Left_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4365__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3327__C _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4668__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3340__A1 net152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Left_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5093__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3643__A2 net363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _1777_ _2208_ _2210_ immu_0.page_table\[13\]\[0\] _2211_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_57_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5780_ _1860_ _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_68_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4731_ _2167_ _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_1172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Left_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4662_ _2057_ _2123_ _2125_ immu_1.page_table\[11\]\[1\] _2127_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6401_ _0783_ clknet_leaf_112_core_clock immu_0.page_table\[15\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3613_ _1308_ net263 _1310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _2069_ _2075_ _2077_ net813 _2085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6332_ _0714_ clknet_leaf_75_core_clock immu_1.page_table\[15\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3544_ net149 net44 _1267_ _1272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_35_core_clock clknet_4_7__leaf_core_clock clknet_leaf_35_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_3_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6263_ _0645_ clknet_leaf_88_core_clock immu_1.page_table\[4\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3475_ _1211_ _1213_ _0895_ _1214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_81_1880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5214_ _1814_ _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_62_1290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6194_ _0576_ clknet_leaf_2_core_clock immu_0.page_table\[11\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5145_ _2269_ _2414_ _2416_ net958 _2420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6649__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5608__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5076_ _2378_ _0107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4027_ _1686_ _1687_ _1416_ _1688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_1050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4831__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input307_I ic0_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6799__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_2082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5978_ _2905_ _0482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3398__A1 _1118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4595__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4929_ _1788_ _2240_ _2284_ _2290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_35_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_74_core_clock clknet_4_11__leaf_core_clock clknet_leaf_74_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5139__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4347__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3428__B _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5311__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3163__B _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output526_I net526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5075__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3625__A2 net269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_1156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5378__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_1419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5109__I _2397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5838__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3260_ _0899_ dmmu1.page_table\[14\]\[4\] _0910_ _1006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3313__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3191_ _0875_ _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6941__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6950_ _0523_ clknet_leaf_56_core_clock dmmu1.page_table\[1\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5901_ _2788_ _2856_ _2858_ dmmu1.page_table\[7\]\[4\] _2863_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_2077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6881_ _0454_ clknet_leaf_67_core_clock dmmu1.page_table\[7\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6015__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ _1796_ _2819_ _2821_ dmmu0.page_table\[1\]\[1\] _2823_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5763_ _2776_ _2778_ _2780_ dmmu1.page_table\[10\]\[0\] _2781_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4714_ _2140_ _2156_ _2158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5447__C _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5694_ _2047_ _2725_ _2727_ net972 _2740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6321__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4329__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4645_ _2116_ _0747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4576_ _2074_ _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5541__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6315_ _0697_ clknet_leaf_70_core_clock dmmu1.page_table\[14\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3527_ net141 net36 _0850_ _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6471__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input257_I dcache_wb_o_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6246_ _0628_ clknet_leaf_84_core_clock immu_1.page_table\[5\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3458_ dmmu1.page_table\[8\]\[10\] dmmu1.page_table\[9\]\[10\] dmmu1.page_table\[10\]\[10\]
+ dmmu1.page_table\[11\]\[10\] _0887_ _0900_ _1198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3304__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4501__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6177_ dmmu1.long_off_reg\[3\] _1852_ _3016_ _3020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3389_ _1129_ _1130_ _0896_ _1131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5128_ _2328_ _2398_ _2400_ immu_0.page_table\[6\]\[8\] _2409_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input20_I c0_o_mem_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5057__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5059_ _2258_ _2367_ _2369_ net812 _2370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4804__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4280__A2 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3466__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3091__I0 net128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3791__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6814__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4335__A3 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7144__I net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6964__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4099__A2 net275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput320 ic0_wb_adr[5] net320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput331 ic1_mem_data[0] net331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3846__A2 _1490_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput342 ic1_mem_data[1] net342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput353 ic1_mem_data[2] net353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold60 dmmu1.page_table\[6\]\[5\] net794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput364 ic1_wb_adr[10] net364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_26_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput375 ic1_wb_adr[6] net375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xhold71 dmmu0.page_table\[8\]\[9\] net805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput386 inner_ext_irq net386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold82 dmmu1.page_table\[9\]\[9\] net816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput397 inner_wb_i_dat[2] net397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_76_1267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold93 dmmu1.page_table\[2\]\[5\] net827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_85_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4271__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6344__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3782__A1 net705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6494__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3209__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4430_ _1985_ _0663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_2 _1262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__A2 _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4361_ _1839_ _1873_ _1892_ _1941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_21_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7054__I net291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6100_ _2974_ _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3312_ dmmu0.page_table\[0\]\[5\] dmmu0.page_table\[1\]\[5\] dmmu0.page_table\[2\]\[5\]
+ dmmu0.page_table\[3\]\[5\] _0864_ _0941_ _1057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_6_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7080_ net333 net486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4292_ _1901_ _0609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5287__A1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6031_ _2849_ _2924_ _2926_ net955 _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3243_ _0932_ _0892_ _0933_ _0989_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_52_1765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3174_ dmmu1.page_table\[8\]\[1\] dmmu1.page_table\[9\]\[1\] dmmu1.page_table\[10\]\[1\]
+ dmmu1.page_table\[11\]\[1\] _0908_ _0910_ _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5039__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6933_ _0506_ clknet_leaf_65_core_clock dmmu1.page_table\[3\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6864_ _0437_ clknet_leaf_51_core_clock dmmu1.page_table\[8\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5815_ _2812_ _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6795_ _0368_ clknet_leaf_47_core_clock dmmu1.page_table\[12\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_2085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _2069_ _2760_ _2762_ dmmu1.page_table\[11\]\[7\] _2770_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4081__C _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5677_ _2731_ _0355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_66_1447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input374_I ic1_wb_adr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4628_ _2105_ _2089_ _2091_ immu_1.page_table\[13\]\[10\] _2106_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6987__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input68_I c0_o_req_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4722__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ _2064_ _0713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_1155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5278__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6229_ _0611_ clknet_leaf_82_core_clock immu_1.page_table\[0\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6367__CLK clknet_leaf_63_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5450__A1 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_2640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_2651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_2662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output593_I net593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7139__I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_1514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5882__I net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_2591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5505__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4308__A3 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_75_2466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3335__C _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__A1 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput150 c1_o_mem_high_addr[0] net150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput161 c1_o_mem_sel[1] net161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput172 c1_o_req_addr[2] net172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3351__B _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput183 c1_sr_bus_addr[11] net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput194 c1_sr_bus_addr[7] net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_1930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_2052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3930_ _1579_ _1582_ _1593_ _1348_ _1594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_54_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3861_ _1375_ _1526_ _1378_ _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7049__I net285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5600_ _2455_ _2681_ _2684_ dmmu0.page_table\[6\]\[3\] _2688_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_45_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6580_ _0153_ clknet_leaf_10_core_clock immu_0.page_table\[4\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5744__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3792_ immu_0.page_table\[4\]\[2\] immu_0.page_table\[5\]\[2\] immu_0.page_table\[6\]\[2\]
+ immu_0.page_table\[7\]\[2\] _1370_ _1372_ _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_15_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5531_ _2300_ _2646_ _2648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4952__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3850__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5462_ _2608_ _0263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_2023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput602 net602 ic0_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_2_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3507__A1 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4413_ net85 net84 _1971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_1_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput613 net613 ic0_wb_i_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__4704__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput624 net624 ic1_mem_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5393_ _2567_ _0235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_58_1963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput635 net635 ic1_mem_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput646 net646 ic1_wb_i_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7132_ net62 net585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4180__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput657 net657 ic1_wb_i_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput668 net668 inner_wb_adr[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4344_ _1932_ _0630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_54_1827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput679 net679 inner_wb_adr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7063_ net301 net452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4275_ _1870_ _1875_ _1877_ immu_1.page_table\[7\]\[10\] _1889_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_35_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6014_ _2927_ _0496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3226_ _0971_ _0972_ _0940_ _0973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_1841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4483__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5680__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3157_ _0906_ _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_input122_I c1_o_mem_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3088_ _0846_ net534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3038__A3 _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5432__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6916_ _0489_ clknet_leaf_56_core_clock dmmu1.page_table\[4\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5983__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6847_ _0420_ clknet_leaf_39_core_clock dmmu0.page_table\[1\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6778_ _0351_ clknet_leaf_104_core_clock dmmu0.long_off_reg\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5729_ _2759_ _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_66_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5408__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5499__A1 _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold360 immu_0.page_table\[10\]\[9\] net1094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold371 dmmu0.page_table\[15\]\[8\] net1105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output439_I net439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_73_core_clock_I clknet_4_9__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5120__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_2047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_2270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_64_2134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_2009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3985__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_2023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3737__A1 net385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_2517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_2539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3832__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6151__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6532__CLK clknet_leaf_6_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4060_ _1368_ _1719_ _1720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4465__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6682__CLK clknet_leaf_100_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4217__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_1620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4962_ _1819_ _2299_ _2302_ dmmu0.page_table\[7\]\[9\] _2312_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_47_1631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5965__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6701_ _0274_ clknet_leaf_35_core_clock dmmu0.page_table\[4\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3913_ net659 net239 _1578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_28_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4893_ _2265_ _2261_ _2263_ dmmu0.page_table\[8\]\[1\] _2266_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_28_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6632_ _0205_ clknet_leaf_33_core_clock dmmu0.page_table\[12\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_15_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5178__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3844_ _1502_ net705 _1505_ _1510_ _1511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_74_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4076__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3728__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6563_ _0136_ clknet_leaf_21_core_clock immu_0.page_table\[5\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3775_ _1433_ _1439_ _1444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_54_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5514_ _2638_ _0285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6494_ _0067_ clknet_leaf_30_core_clock dmmu0.page_table\[14\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5445_ _2597_ _0257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput410 net410 c0_i_mem_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput421 net421 c0_i_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_30_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput432 net432 c0_i_req_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput443 net443 c0_i_req_data[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4153__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5350__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5376_ _2455_ _2553_ _2555_ net890 _2559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput454 net454 c0_i_req_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput465 net465 c1_i_mc_core_int vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput476 net476 c1_i_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7115_ net391 net568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput487 net487 c1_i_req_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4327_ _1864_ _1911_ _1914_ net975 _1922_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput498 net498 c1_i_req_data[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3770__I _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input337_I ic1_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7046_ net282 net433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4258_ _1880_ _0596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_38_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3209_ dmmu0.page_table\[0\]\[2\] dmmu0.page_table\[1\]\[2\] dmmu0.page_table\[2\]\[2\]
+ dmmu0.page_table\[3\]\[2\] _0950_ _0952_ _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4189_ _1823_ _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_69_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3211__S _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3967__A1 net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_2007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5708__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3719__A1 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6555__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold190 dmmu1.page_table\[13\]\[1\] net924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_79_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7152__I net392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5644__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Right_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_1143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3502__S0 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3186__A2 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4383__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3560_ net161 net56 _0841_ _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_25_Right_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_25_core_clock clknet_4_5__leaf_core_clock clknet_leaf_25_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3491_ net51 dmmu0.long_off_reg\[6\] _1229_ _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_23_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5230_ _2451_ _2470_ _2472_ immu_0.page_table\[2\]\[1\] _2474_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_36_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5883__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5161_ _1972_ _2296_ _2428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_20_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4112_ _1765_ _1766_ _1767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5092_ _2388_ _0113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4043_ immu_0.page_table\[0\]\[9\] immu_0.page_table\[1\]\[9\] immu_0.page_table\[2\]\[9\]
+ immu_0.page_table\[3\]\[9\] _1396_ _1371_ _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_79_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Right_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3741__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6428__CLK clknet_leaf_110_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5994_ _2915_ _0488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_1063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4945_ _2303_ _0051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_23_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4876_ _1819_ _2242_ _2244_ net852 _2254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_64_core_clock clknet_4_11__leaf_core_clock clknet_leaf_64_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6578__CLK clknet_leaf_24_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3827_ _1463_ immu_0.page_table\[15\]\[3\] _1494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6615_ _0188_ clknet_leaf_8_core_clock immu_0.page_table\[0\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3765__I _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Right_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5410__I1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3177__A2 _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input287_I ic0_mem_data[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6546_ _0119_ clknet_leaf_21_core_clock immu_0.page_table\[7\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_2084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3758_ _1382_ _1426_ _1372_ _1427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__5571__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6477_ _0050_ clknet_leaf_105_core_clock net407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_42_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5980__I _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6115__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3689_ _1350_ net310 _1360_ _1361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4126__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5428_ _2457_ _2582_ _2584_ dmmu0.page_table\[2\]\[4\] _2589_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input50_I c0_o_mem_high_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5874__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5359_ _2548_ _0220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3206__S _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Right_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5626__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4429__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7029_ net384 net405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_69_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5929__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_2004 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4601__A2 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_2000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3675__I _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7147__I net402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4365__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_1309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4668__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_70_Right_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5093__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6720__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5396__A3 _1971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4730_ _1815_ _2157_ _2159_ net965 _2167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_57_966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4661_ _2126_ _0753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6400_ _0782_ clknet_leaf_111_core_clock immu_0.page_table\[15\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3612_ _1309_ net685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6870__CLK clknet_leaf_68_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4592_ _2084_ _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6331_ _0713_ clknet_leaf_77_core_clock immu_1.page_table\[15\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3543_ _1271_ net557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6262_ _0644_ clknet_leaf_87_core_clock immu_1.page_table\[4\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3474_ _0906_ _1212_ _0912_ _1213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5856__A1 _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5213_ _2462_ _0160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6193_ _0575_ clknet_leaf_9_core_clock immu_0.page_table\[11\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5144_ _2419_ _0134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3253__C _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5608__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5459__I1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6250__CLK clknet_leaf_85_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5075_ _2328_ _2367_ _2369_ net956 _2378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4026_ immu_1.page_table\[4\]\[9\] immu_1.page_table\[5\]\[9\] immu_1.page_table\[6\]\[9\]
+ immu_1.page_table\[7\]\[9\] _1441_ _1442_ _1687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_79_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4831__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input202_I c1_sr_bus_data_o[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6033__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ net200 _2889_ _2891_ net1070 _2905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4595__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3398__A2 _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4928_ net406 _2288_ _2289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input98_I c0_sr_bus_data_o[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3709__B _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4859_ _2245_ _0023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4347__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6529_ _0102_ clknet_leaf_9_core_clock immu_0.page_table\[8\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_2010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_12_core_clock_I clknet_4_3__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3444__B _1119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3173__I2 dmmu1.page_table\[14\]\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6743__CLK clknet_leaf_42_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3228__I3 dmmu0.page_table\[7\]\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6893__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5535__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5838__A1 _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6273__CLK clknet_leaf_90_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3190_ _0936_ _0937_ _0938_ _0939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5900_ _2862_ _0447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6880_ _0453_ clknet_leaf_59_core_clock dmmu1.page_table\[7\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6015__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ _2822_ _0418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4577__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5762_ _2779_ _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_72_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4713_ _2156_ _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_17_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5693_ _2739_ _0363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_1965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4329__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4204__I _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4644_ _2065_ _2108_ _2110_ immu_1.page_table\[12\]\[5\] _2116_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3248__C _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4575_ _1838_ _1909_ _2028_ _2074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_12_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6616__CLK clknet_leaf_17_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3526_ _1262_ net543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6314_ _0696_ clknet_leaf_70_core_clock dmmu1.page_table\[14\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_core_clock_I clknet_4_1__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6245_ _0627_ clknet_leaf_94_core_clock immu_1.page_table\[2\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3457_ _0896_ _1196_ _1197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_111_core_clock clknet_4_0__leaf_core_clock clknet_leaf_111_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input152_I c1_o_mem_high_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4501__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6176_ _3019_ _0566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3388_ dmmu1.page_table\[4\]\[8\] dmmu1.page_table\[5\]\[8\] dmmu1.page_table\[6\]\[8\]
+ dmmu1.page_table\[7\]\[8\] _0898_ _0909_ _1130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5127_ _2408_ _0128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_1736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_78_core_clock_I clknet_4_11__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_2_Right_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3068__A1 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5058_ _2368_ _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_58_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input13_I c0_o_mem_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4265__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4804__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4009_ immu_0.page_table\[0\]\[8\] immu_0.page_table\[1\]\[8\] immu_0.page_table\[2\]\[8\]
+ immu_0.page_table\[3\]\[8\] _1487_ _1455_ _1671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_32_2009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A3 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4032__A3 _1692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3091__I1 net23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4114__I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5517__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_1562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_73_Left_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_2394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3926__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput310 ic0_wb_adr[10] net310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_60_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput321 ic0_wb_adr[6] net321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3846__A3 _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput332 ic1_mem_data[10] net332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput343 ic1_mem_data[20] net343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput354 ic1_mem_data[30] net354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_1213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold50 dmmu1.page_table\[1\]\[2\] net784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__7160__I net174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput365 ic1_wb_adr[11] net365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput376 ic1_wb_adr[7] net376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold61 immu_1.page_table\[15\]\[1\] net795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_56_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold72 dmmu0.page_table\[10\]\[12\] net806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold83 dmmu1.page_table\[6\]\[6\] net817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput387 inner_wb_ack net387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3059__A1 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput398 inner_wb_i_dat[3] net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xhold94 dmmu1.page_table\[2\]\[12\] net828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_19_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_82_Left_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_80_core_clock_I clknet_4_10__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3231__A1 _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6639__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_3 _1276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4360_ _1940_ _0638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6789__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3311_ _0940_ _1055_ _0879_ _1056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4291_ _1851_ _1894_ _1897_ immu_1.page_table\[0\]\[3\] _1901_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_24_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6030_ _2935_ _0504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5287__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3242_ _0974_ _0979_ _0984_ _0988_ net523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_TAPCELL_ROW_56_1891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I c0_o_instr_long_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4495__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3173_ dmmu1.page_table\[12\]\[1\] dmmu1.page_table\[13\]\[1\] dmmu1.page_table\[14\]\[1\]
+ dmmu1.page_table\[15\]\[1\] _0908_ _0902_ _0922_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_52_1777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5039__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4798__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6932_ _0505_ clknet_leaf_62_core_clock dmmu1.page_table\[3\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3103__I _0854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5995__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6863_ _0436_ clknet_leaf_51_core_clock dmmu1.page_table\[8\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3470__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5814_ _2794_ _2802_ _2804_ net830 _2812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6794_ _0367_ clknet_leaf_47_core_clock dmmu1.page_table\[12\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5745_ _2769_ _0385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3222__A1 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5676_ _2059_ _2726_ _2728_ net1052 _2731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4627_ net198 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3773__I _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4722__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input367_I ic1_wb_adr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4558_ _2063_ _2053_ _2055_ net739 _2064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3509_ net156 dmmu1.long_off_reg\[6\] _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4489_ _1852_ _2014_ _2016_ immu_1.page_table\[3\]\[3\] _2020_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _0610_ clknet_leaf_84_core_clock immu_1.page_table\[0\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3722__B _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6159_ _1863_ _3000_ _3002_ net1031 _3010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_55_1831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5450__A2 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_2641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3300__I2 dmmu1.page_table\[14\]\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3461__A1 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_2652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_2663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5738__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3213__A1 _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output586_I net586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_11_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6163__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7155__I net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_2456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5269__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput140 c1_o_mem_data[15] net140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput151 c1_o_mem_high_addr[1] net151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput162 c1_o_mem_we net162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput173 c1_o_req_addr[3] net173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6311__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput184 c1_sr_bus_addr[12] net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput195 c1_sr_bus_addr[8] net195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4229__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6461__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3860_ immu_0.page_table\[4\]\[4\] immu_0.page_table\[5\]\[4\] immu_0.page_table\[6\]\[4\]
+ immu_0.page_table\[7\]\[4\] _1396_ _1371_ _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_58_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_12__f_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3791_ _1382_ _1458_ _1375_ _1459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_45_1581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4401__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4952__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5530_ _2646_ _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_41_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5461_ immu_1.high_addr_off\[4\] _1855_ _2603_ _2608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7065__I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4412_ _1970_ _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput603 net603 ic0_wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__4704__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput614 net614 ic0_wb_i_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5392_ _1994_ _2552_ _2554_ net846 _2567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5901__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput625 net625 ic1_mem_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput636 net636 ic1_mem_cache_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput647 net647 ic1_wb_i_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7131_ net61 net584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4343_ _1849_ _1927_ _1929_ immu_1.page_table\[5\]\[2\] _1932_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput658 net658 inner_wb_4_burst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4180__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput669 net669 inner_wb_adr[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7062_ net300 net451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4274_ _1888_ _0604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6013_ _2776_ _2924_ _2926_ dmmu1.page_table\[3\]\[0\] _2927_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3225_ dmmu0.page_table\[12\]\[3\] dmmu0.page_table\[13\]\[3\] dmmu0.page_table\[14\]\[3\]
+ dmmu0.page_table\[15\]\[3\] _0950_ _0952_ _0972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_20_1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5680__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3156_ _0905_ _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3087_ net126 net21 _0842_ _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6804__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input115_I c1_o_instr_long_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5432__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6915_ _0488_ clknet_leaf_57_core_clock dmmu1.page_table\[4\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4640__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6846_ _0419_ clknet_leaf_43_core_clock dmmu0.page_table\[1\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6777_ _0350_ clknet_leaf_103_core_clock dmmu0.long_off_reg\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3989_ _1616_ _1649_ _1650_ _1651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_45_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5728_ _1826_ _1874_ _2031_ _2759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA_input80_I c0_sr_bus_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6145__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5659_ _2720_ _0348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold350 immu_1.page_table\[11\]\[5\] net1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold361 immu_0.page_table\[5\]\[8\] net1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold372 immu_0.page_table\[10\]\[8\] net1106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6334__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4459__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5120__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_5_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output501_I net501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_2714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6484__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5959__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_2271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_64_2146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3985__A2 net241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4934__A1 net407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_2518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_core_clock clknet_4_6__leaf_core_clock clknet_leaf_15_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_2074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4870__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6977__CLK clknet_leaf_105_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4961_ _2311_ _0059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3425__A1 _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4622__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ _0273_ clknet_leaf_41_core_clock dmmu0.page_table\[4\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3912_ _1552_ _1576_ _1577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_1133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_28_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4892_ _1796_ _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_54_core_clock clknet_4_15__leaf_core_clock clknet_leaf_54_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_28_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6631_ _0204_ clknet_leaf_38_core_clock dmmu0.page_table\[12\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5178__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3843_ _1433_ _1506_ _1509_ _1434_ _1510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_46_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6207__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3774_ immu_1.page_table\[4\]\[1\] immu_1.page_table\[5\]\[1\] immu_1.page_table\[6\]\[1\]
+ immu_1.page_table\[7\]\[1\] _1441_ _1442_ _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_27_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6562_ _0135_ clknet_leaf_27_core_clock immu_0.page_table\[5\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5513_ _2459_ _2630_ _2632_ net997 _2638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6493_ _0066_ clknet_leaf_30_core_clock dmmu0.page_table\[14\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4212__I _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5444_ _1996_ _2581_ _2583_ dmmu0.page_table\[2\]\[12\] _2597_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput411 net411 c0_i_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6357__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput422 net422 c0_i_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput433 net433 c0_i_req_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5350__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput444 net444 c0_i_req_data[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4153__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput455 net455 c0_i_req_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5375_ _2558_ _0226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput466 net466 c1_i_mem_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7114_ net390 net567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput477 net477 c1_i_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput488 net488 c1_i_req_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4326_ _1921_ _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput499 net499 c1_i_req_data[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_leaf_17_core_clock_I clknet_4_5__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4257_ _1846_ _1876_ _1878_ net1080 _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7045_ net281 net432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input232_I dcache_wb_adr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3208_ dmmu0.page_table\[8\]\[2\] dmmu0.page_table\[9\]\[2\] dmmu0.page_table\[10\]\[2\]
+ dmmu0.page_table\[11\]\[2\] _0950_ _0952_ _0956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_39_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4188_ net197 _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_1683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3139_ _0888_ _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_1547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4613__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6829_ _0402_ clknet_leaf_69_core_clock dmmu1.page_table\[10\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_1529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6133__A3 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output451_I net451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_2085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold180 dmmu0.page_table\[9\]\[3\] net914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold191 dmmu0.page_table\[12\]\[0\] net925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5644__A2 _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_2208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_2023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3502__S1 net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4080__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6109__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4383__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3490_ _1180_ _1183_ _1228_ _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_80_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_1197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5332__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_36_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5160_ _2427_ _0142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_8_core_clock_I clknet_4_1__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4111_ icache_arbiter.o_sel_sig net379 _1766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5091_ _2269_ _2382_ _2384_ net797 _2388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4042_ immu_0.page_table\[4\]\[9\] immu_0.page_table\[5\]\[9\] immu_0.page_table\[6\]\[9\]
+ immu_0.page_table\[7\]\[9\] _1396_ _1371_ _1703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__3646__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4843__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3741__S1 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5993_ _2790_ _2907_ _2909_ dmmu1.page_table\[4\]\[5\] _2915_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _2258_ _2299_ _2302_ dmmu0.page_table\[7\]\[0\] _2303_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_23_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4875_ _2253_ _0031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6614_ _0187_ clknet_leaf_20_core_clock immu_0.page_table\[0\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3826_ _1385_ immu_0.page_table\[14\]\[3\] _1493_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_1649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6545_ _0118_ clknet_leaf_23_core_clock immu_0.page_table\[7\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5571__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3757_ _1423_ _1425_ _1366_ _1426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input182_I c1_sr_bus_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6476_ _0049_ clknet_leaf_92_core_clock net406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_3688_ _1304_ _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_28_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4126__A2 _0815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5427_ _2588_ _0248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_7_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5874__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4098__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5358_ _2529_ _2536_ _2538_ dmmu0.page_table\[15\]\[9\] _2548_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input43_I c0_o_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4309_ _1910_ _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5087__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5289_ _1805_ _2502_ _2504_ immu_0.page_table\[0\]\[4\] _2508_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5626__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3637__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6051__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4062__A1 _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4601__A3 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6522__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output499_I net499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5011__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_2001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_85_core_clock_I clknet_4_10__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4365__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6672__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7163__I net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3420__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_17_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3100__I0 net132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5396__A4 _1972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_5_core_clock clknet_4_1__leaf_core_clock clknet_leaf_5_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3800__A1 _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4660_ _2051_ _2123_ _2125_ net927 _2126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3239__S0 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3611_ _1308_ net256 _1309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5553__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4591_ _2067_ _2075_ _2077_ net978 _2084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _0712_ clknet_leaf_72_core_clock immu_1.page_table\[15\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3542_ net148 net43 _1267_ _1271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1092 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5305__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6261_ _0643_ clknet_leaf_85_core_clock immu_1.page_table\[4\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3473_ dmmu1.page_table\[0\]\[11\] dmmu1.page_table\[1\]\[11\] dmmu1.page_table\[2\]\[11\]
+ dmmu1.page_table\[3\]\[11\] _0898_ _0901_ _1212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__7073__I net357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_101_core_clock clknet_4_2__leaf_core_clock clknet_leaf_101_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_23_1210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5856__A2 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5212_ _2461_ _2447_ _2449_ immu_0.page_table\[3\]\[6\] _2462_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3867__A1 net5 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6192_ _0574_ clknet_leaf_7_core_clock immu_0.page_table\[11\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5143_ _2267_ _2414_ _2416_ immu_0.page_table\[5\]\[2\] _2419_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5069__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5608__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5074_ _2377_ _0106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3619__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4816__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4025_ immu_1.page_table\[0\]\[9\] immu_1.page_table\[1\]\[9\] immu_1.page_table\[2\]\[9\]
+ immu_1.page_table\[3\]\[9\] _1441_ _1442_ _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_56_1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__CLK clknet_leaf_23_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6033__A2 _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5976_ _2904_ _0481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4927_ _1776_ _2285_ _2287_ _1823_ _2288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4595__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5792__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input397_I inner_wb_i_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4858_ _1777_ _2242_ _2244_ net1017 _2245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4347__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3809_ immu_1.page_table\[12\]\[2\] immu_1.page_table\[13\]\[2\] _1474_ _1477_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4789_ _2202_ _0805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6528_ _0101_ clknet_leaf_7_core_clock immu_0.page_table\[8\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3725__B _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6459_ _0032_ clknet_leaf_12_core_clock dmmu0.page_table\[9\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_2044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4283__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4035__A1 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5232__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7158__I net172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5535__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__CLK clknet_leaf_109_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5299__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4310__I _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5838__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_2095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_2057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6015__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6173__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5830_ _1776_ _2819_ _2821_ dmmu0.page_table\[1\]\[0\] _2822_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5761_ _2682_ _2777_ _2779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7068__I net407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ _1790_ _2155_ _2156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_31_1556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5692_ _2105_ _2725_ _2727_ dmmu1.page_table\[13\]\[10\] _2739_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4329__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4643_ _2115_ _0746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4574_ _2073_ _0719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6313_ _0695_ clknet_leaf_94_core_clock immu_1.page_table\[3\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3525_ net134 net29 _0850_ _1262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4220__I _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6244_ _0626_ clknet_leaf_88_core_clock immu_1.page_table\[2\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3264__C _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3456_ dmmu1.page_table\[12\]\[10\] dmmu1.page_table\[13\]\[10\] dmmu1.page_table\[14\]\[10\]
+ dmmu1.page_table\[15\]\[10\] _0887_ _0900_ _1196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_42_1652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4501__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6175_ dmmu1.long_off_reg\[2\] _1849_ _3016_ _3019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3387_ dmmu1.page_table\[0\]\[8\] dmmu1.page_table\[1\]\[8\] dmmu1.page_table\[2\]\[8\]
+ dmmu1.page_table\[3\]\[8\] _0898_ _0909_ _1129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3560__I0 net161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input145_I c1_o_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5126_ _2277_ _2398_ _2400_ immu_0.page_table\[6\]\[7\] _2408_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5057_ _2140_ _2366_ _2368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3068__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4265__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input312_I ic0_wb_adr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4008_ immu_0.page_table\[4\]\[8\] immu_0.page_table\[5\]\[8\] immu_0.page_table\[6\]\[8\]
+ immu_0.page_table\[7\]\[8\] _1424_ _1455_ _1670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_71_1325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4017__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5959_ _2786_ _2890_ _2892_ dmmu1.page_table\[5\]\[3\] _2896_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3439__C _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5517__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6710__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_2395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output629_I net629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput300 ic0_mem_data[30] net300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3926__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput311 ic0_wb_adr[11] net311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput322 ic0_wb_adr[7] net322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput333 ic1_mem_data[11] net333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput344 ic1_mem_data[21] net344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold40 dmmu1.page_table\[6\]\[10\] net774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput355 ic1_mem_data[31] net355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold51 immu_1.page_table\[8\]\[9\] net785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold62 dmmu1.page_table\[1\]\[11\] net796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput366 ic1_wb_adr[12] net366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput377 ic1_wb_adr[8] net377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold73 dmmu1.page_table\[3\]\[12\] net807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput388 inner_wb_err net388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput399 inner_wb_i_dat[4] net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3059__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold84 immu_0.page_table\[6\]\[10\] net818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6860__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold95 immu_1.page_table\[10\]\[9\] net829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_54_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5756__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3349__C _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3231__A2 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3862__S0 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6240__CLK clknet_leaf_89_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_4 net373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3310_ dmmu0.page_table\[8\]\[5\] dmmu0.page_table\[9\]\[5\] dmmu0.page_table\[10\]\[5\]
+ dmmu0.page_table\[11\]\[5\] _0865_ _0868_ _1055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_4290_ _1900_ _0608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3241_ _0895_ _0987_ _0915_ _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_1972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4495__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3542__I0 net148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3172_ _0881_ _0885_ _0921_ _0822_ net520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_TAPCELL_ROW_52_1767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5444__B1 _2583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6931_ _0504_ clknet_leaf_60_core_clock dmmu1.page_table\[3\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5995__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4798__A2 _2207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _0435_ clknet_leaf_50_core_clock dmmu1.page_table\[8\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5813_ _2811_ _0411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6793_ _0366_ clknet_leaf_47_core_clock dmmu1.page_table\[12\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5744_ _2067_ _2760_ _2762_ dmmu1.page_table\[11\]\[6\] _2769_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3853__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5675_ _2730_ _0354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4626_ _2104_ _0740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_83_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6733__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4722__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4557_ _1854_ _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_64_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input262_I dcache_wb_o_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3508_ _1119_ _1236_ _1245_ _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4488_ _2019_ _0687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6227_ _0609_ clknet_leaf_90_core_clock immu_1.page_table\[0\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3439_ _0878_ _1173_ _1178_ _0862_ _1179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_42_1471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4030__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6883__CLK clknet_leaf_68_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3533__I0 net144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6158_ _3009_ _0558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5109_ _2397_ _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_38_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6089_ _2847_ _2958_ _2960_ dmmu1.page_table\[1\]\[8\] _2969_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3230__S _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_2642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3461__A2 _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_2653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5738__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6263__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_24_core_clock_I clknet_4_5__leaf_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6163__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_2479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7171__I net170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4477__A1 net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5674__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput130 c1_o_mem_addr[6] net130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput141 c1_o_mem_data[1] net141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput152 c1_o_mem_high_addr[2] net152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput163 c1_o_req_active net163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_21_1588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput174 c1_o_req_addr[4] net174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4229__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3204__I _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput185 c1_sr_bus_addr[13] net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5426__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput196 c1_sr_bus_addr[9] net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5977__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6606__CLK clknet_leaf_24_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_44_core_clock clknet_4_12__leaf_core_clock clknet_leaf_44_core_clock
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_85_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4401__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3790_ _1456_ _1457_ _1377_ _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6756__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4952__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5460_ _2607_ _0262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_2101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4411_ _1870_ _1956_ _1958_ immu_1.page_table\[6\]\[10\] _1970_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4165__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput604 net604 ic0_wb_i_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4704__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5901__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _2566_ _0234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput615 net615 ic0_wb_i_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_58_1954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput626 net626 ic1_mem_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput637 net637 ic1_mem_ppl_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7130_ net60 net583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_58_1965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4342_ _1931_ _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput648 net648 ic1_wb_i_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput659 net659 inner_wb_8_burst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3823__B _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7061_ net298 net449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_39_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4273_ _1868_ _1876_ _1878_ immu_1.page_table\[7\]\[9\] _1888_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7081__I net334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6012_ _2925_ _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3224_ dmmu0.page_table\[8\]\[3\] dmmu0.page_table\[9\]\[3\] dmmu0.page_table\[10\]\[3\]
+ dmmu0.page_table\[11\]\[3\] _0950_ _0948_ _0971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
.ends

