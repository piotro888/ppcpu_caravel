magic
tech sky130B
magscale 1 2
timestamp 1663070888
<< nwell >>
rect 1066 37253 38862 37574
rect 1066 36165 38862 36731
rect 1066 35077 38862 35643
rect 1066 33989 38862 34555
rect 1066 32901 38862 33467
rect 1066 31813 38862 32379
rect 1066 30725 38862 31291
rect 1066 29637 38862 30203
rect 1066 28549 38862 29115
rect 1066 27461 38862 28027
rect 1066 26373 38862 26939
rect 1066 25285 38862 25851
rect 1066 24197 38862 24763
rect 1066 23109 38862 23675
rect 1066 22021 38862 22587
rect 1066 20933 38862 21499
rect 1066 19845 38862 20411
rect 1066 18757 38862 19323
rect 1066 17669 38862 18235
rect 1066 16581 38862 17147
rect 1066 15493 38862 16059
rect 1066 14405 38862 14971
rect 1066 13317 38862 13883
rect 1066 12229 38862 12795
rect 1066 11141 38862 11707
rect 1066 10053 38862 10619
rect 1066 8965 38862 9531
rect 1066 7877 38862 8443
rect 1066 6789 38862 7355
rect 1066 5701 38862 6267
rect 1066 4613 38862 5179
rect 1066 3525 38862 4091
rect 1066 2437 38862 3003
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 1104 2128 38824 37584
<< metal2 >>
rect 2318 39200 2374 40000
rect 3054 39200 3110 40000
rect 3790 39200 3846 40000
rect 4526 39200 4582 40000
rect 5262 39200 5318 40000
rect 5998 39200 6054 40000
rect 6734 39200 6790 40000
rect 7470 39200 7526 40000
rect 8206 39200 8262 40000
rect 8942 39200 8998 40000
rect 9678 39200 9734 40000
rect 10414 39200 10470 40000
rect 11150 39200 11206 40000
rect 11886 39200 11942 40000
rect 12622 39200 12678 40000
rect 13358 39200 13414 40000
rect 14094 39200 14150 40000
rect 14830 39200 14886 40000
rect 15566 39200 15622 40000
rect 16302 39200 16358 40000
rect 17038 39200 17094 40000
rect 17774 39200 17830 40000
rect 18510 39200 18566 40000
rect 19246 39200 19302 40000
rect 19982 39200 20038 40000
rect 20718 39200 20774 40000
rect 21454 39200 21510 40000
rect 22190 39200 22246 40000
rect 22926 39200 22982 40000
rect 23662 39200 23718 40000
rect 24398 39200 24454 40000
rect 25134 39200 25190 40000
rect 25870 39200 25926 40000
rect 26606 39200 26662 40000
rect 27342 39200 27398 40000
rect 28078 39200 28134 40000
rect 28814 39200 28870 40000
rect 29550 39200 29606 40000
rect 30286 39200 30342 40000
rect 31022 39200 31078 40000
rect 31758 39200 31814 40000
rect 32494 39200 32550 40000
rect 33230 39200 33286 40000
rect 33966 39200 34022 40000
rect 34702 39200 34758 40000
rect 35438 39200 35494 40000
rect 36174 39200 36230 40000
rect 36910 39200 36966 40000
rect 37646 39200 37702 40000
rect 2318 0 2374 800
rect 3054 0 3110 800
rect 3790 0 3846 800
rect 4526 0 4582 800
rect 5262 0 5318 800
rect 5998 0 6054 800
rect 6734 0 6790 800
rect 7470 0 7526 800
rect 8206 0 8262 800
rect 8942 0 8998 800
rect 9678 0 9734 800
rect 10414 0 10470 800
rect 11150 0 11206 800
rect 11886 0 11942 800
rect 12622 0 12678 800
rect 13358 0 13414 800
rect 14094 0 14150 800
rect 14830 0 14886 800
rect 15566 0 15622 800
rect 16302 0 16358 800
rect 17038 0 17094 800
rect 17774 0 17830 800
rect 18510 0 18566 800
rect 19246 0 19302 800
rect 19982 0 20038 800
rect 20718 0 20774 800
rect 21454 0 21510 800
rect 22190 0 22246 800
rect 22926 0 22982 800
rect 23662 0 23718 800
rect 24398 0 24454 800
rect 25134 0 25190 800
rect 25870 0 25926 800
rect 26606 0 26662 800
rect 27342 0 27398 800
rect 28078 0 28134 800
rect 28814 0 28870 800
rect 29550 0 29606 800
rect 30286 0 30342 800
rect 31022 0 31078 800
rect 31758 0 31814 800
rect 32494 0 32550 800
rect 33230 0 33286 800
rect 33966 0 34022 800
rect 34702 0 34758 800
rect 35438 0 35494 800
rect 36174 0 36230 800
rect 36910 0 36966 800
rect 37646 0 37702 800
<< obsm2 >>
rect 2430 39144 2998 39250
rect 3166 39144 3734 39250
rect 3902 39144 4470 39250
rect 4638 39144 5206 39250
rect 5374 39144 5942 39250
rect 6110 39144 6678 39250
rect 6846 39144 7414 39250
rect 7582 39144 8150 39250
rect 8318 39144 8886 39250
rect 9054 39144 9622 39250
rect 9790 39144 10358 39250
rect 10526 39144 11094 39250
rect 11262 39144 11830 39250
rect 11998 39144 12566 39250
rect 12734 39144 13302 39250
rect 13470 39144 14038 39250
rect 14206 39144 14774 39250
rect 14942 39144 15510 39250
rect 15678 39144 16246 39250
rect 16414 39144 16982 39250
rect 17150 39144 17718 39250
rect 17886 39144 18454 39250
rect 18622 39144 19190 39250
rect 19358 39144 19926 39250
rect 20094 39144 20662 39250
rect 20830 39144 21398 39250
rect 21566 39144 22134 39250
rect 22302 39144 22870 39250
rect 23038 39144 23606 39250
rect 23774 39144 24342 39250
rect 24510 39144 25078 39250
rect 25246 39144 25814 39250
rect 25982 39144 26550 39250
rect 26718 39144 27286 39250
rect 27454 39144 28022 39250
rect 28190 39144 28758 39250
rect 28926 39144 29494 39250
rect 29662 39144 30230 39250
rect 30398 39144 30966 39250
rect 31134 39144 31702 39250
rect 31870 39144 32438 39250
rect 32606 39144 33174 39250
rect 33342 39144 33910 39250
rect 34078 39144 34646 39250
rect 34814 39144 35382 39250
rect 35550 39144 36118 39250
rect 36286 39144 36854 39250
rect 37022 39144 37590 39250
rect 37758 39144 38252 39250
rect 2320 856 38252 39144
rect 2430 800 2998 856
rect 3166 800 3734 856
rect 3902 800 4470 856
rect 4638 800 5206 856
rect 5374 800 5942 856
rect 6110 800 6678 856
rect 6846 800 7414 856
rect 7582 800 8150 856
rect 8318 800 8886 856
rect 9054 800 9622 856
rect 9790 800 10358 856
rect 10526 800 11094 856
rect 11262 800 11830 856
rect 11998 800 12566 856
rect 12734 800 13302 856
rect 13470 800 14038 856
rect 14206 800 14774 856
rect 14942 800 15510 856
rect 15678 800 16246 856
rect 16414 800 16982 856
rect 17150 800 17718 856
rect 17886 800 18454 856
rect 18622 800 19190 856
rect 19358 800 19926 856
rect 20094 800 20662 856
rect 20830 800 21398 856
rect 21566 800 22134 856
rect 22302 800 22870 856
rect 23038 800 23606 856
rect 23774 800 24342 856
rect 24510 800 25078 856
rect 25246 800 25814 856
rect 25982 800 26550 856
rect 26718 800 27286 856
rect 27454 800 28022 856
rect 28190 800 28758 856
rect 28926 800 29494 856
rect 29662 800 30230 856
rect 30398 800 30966 856
rect 31134 800 31702 856
rect 31870 800 32438 856
rect 32606 800 33174 856
rect 33342 800 33910 856
rect 34078 800 34646 856
rect 34814 800 35382 856
rect 35550 800 36118 856
rect 36286 800 36854 856
rect 37022 800 37590 856
rect 37758 800 38252 856
<< metal3 >>
rect 39200 37272 40000 37392
rect 39200 36592 40000 36712
rect 39200 35912 40000 36032
rect 39200 35232 40000 35352
rect 39200 34552 40000 34672
rect 39200 33872 40000 33992
rect 39200 33192 40000 33312
rect 39200 32512 40000 32632
rect 39200 31832 40000 31952
rect 39200 31152 40000 31272
rect 39200 30472 40000 30592
rect 39200 29792 40000 29912
rect 39200 29112 40000 29232
rect 39200 28432 40000 28552
rect 39200 27752 40000 27872
rect 39200 27072 40000 27192
rect 39200 26392 40000 26512
rect 39200 25712 40000 25832
rect 39200 25032 40000 25152
rect 39200 24352 40000 24472
rect 39200 23672 40000 23792
rect 39200 22992 40000 23112
rect 39200 22312 40000 22432
rect 39200 21632 40000 21752
rect 39200 20952 40000 21072
rect 39200 20272 40000 20392
rect 39200 19592 40000 19712
rect 39200 18912 40000 19032
rect 39200 18232 40000 18352
rect 39200 17552 40000 17672
rect 39200 16872 40000 16992
rect 39200 16192 40000 16312
rect 39200 15512 40000 15632
rect 39200 14832 40000 14952
rect 39200 14152 40000 14272
rect 39200 13472 40000 13592
rect 39200 12792 40000 12912
rect 39200 12112 40000 12232
rect 39200 11432 40000 11552
rect 39200 10752 40000 10872
rect 39200 10072 40000 10192
rect 39200 9392 40000 9512
rect 39200 8712 40000 8832
rect 39200 8032 40000 8152
rect 39200 7352 40000 7472
rect 39200 6672 40000 6792
rect 39200 5992 40000 6112
rect 39200 5312 40000 5432
rect 39200 4632 40000 4752
rect 39200 3952 40000 4072
rect 39200 3272 40000 3392
rect 39200 2592 40000 2712
<< obsm3 >>
rect 4210 37472 39200 37569
rect 4210 37192 39120 37472
rect 4210 36792 39200 37192
rect 4210 36512 39120 36792
rect 4210 36112 39200 36512
rect 4210 35832 39120 36112
rect 4210 35432 39200 35832
rect 4210 35152 39120 35432
rect 4210 34752 39200 35152
rect 4210 34472 39120 34752
rect 4210 34072 39200 34472
rect 4210 33792 39120 34072
rect 4210 33392 39200 33792
rect 4210 33112 39120 33392
rect 4210 32712 39200 33112
rect 4210 32432 39120 32712
rect 4210 32032 39200 32432
rect 4210 31752 39120 32032
rect 4210 31352 39200 31752
rect 4210 31072 39120 31352
rect 4210 30672 39200 31072
rect 4210 30392 39120 30672
rect 4210 29992 39200 30392
rect 4210 29712 39120 29992
rect 4210 29312 39200 29712
rect 4210 29032 39120 29312
rect 4210 28632 39200 29032
rect 4210 28352 39120 28632
rect 4210 27952 39200 28352
rect 4210 27672 39120 27952
rect 4210 27272 39200 27672
rect 4210 26992 39120 27272
rect 4210 26592 39200 26992
rect 4210 26312 39120 26592
rect 4210 25912 39200 26312
rect 4210 25632 39120 25912
rect 4210 25232 39200 25632
rect 4210 24952 39120 25232
rect 4210 24552 39200 24952
rect 4210 24272 39120 24552
rect 4210 23872 39200 24272
rect 4210 23592 39120 23872
rect 4210 23192 39200 23592
rect 4210 22912 39120 23192
rect 4210 22512 39200 22912
rect 4210 22232 39120 22512
rect 4210 21832 39200 22232
rect 4210 21552 39120 21832
rect 4210 21152 39200 21552
rect 4210 20872 39120 21152
rect 4210 20472 39200 20872
rect 4210 20192 39120 20472
rect 4210 19792 39200 20192
rect 4210 19512 39120 19792
rect 4210 19112 39200 19512
rect 4210 18832 39120 19112
rect 4210 18432 39200 18832
rect 4210 18152 39120 18432
rect 4210 17752 39200 18152
rect 4210 17472 39120 17752
rect 4210 17072 39200 17472
rect 4210 16792 39120 17072
rect 4210 16392 39200 16792
rect 4210 16112 39120 16392
rect 4210 15712 39200 16112
rect 4210 15432 39120 15712
rect 4210 15032 39200 15432
rect 4210 14752 39120 15032
rect 4210 14352 39200 14752
rect 4210 14072 39120 14352
rect 4210 13672 39200 14072
rect 4210 13392 39120 13672
rect 4210 12992 39200 13392
rect 4210 12712 39120 12992
rect 4210 12312 39200 12712
rect 4210 12032 39120 12312
rect 4210 11632 39200 12032
rect 4210 11352 39120 11632
rect 4210 10952 39200 11352
rect 4210 10672 39120 10952
rect 4210 10272 39200 10672
rect 4210 9992 39120 10272
rect 4210 9592 39200 9992
rect 4210 9312 39120 9592
rect 4210 8912 39200 9312
rect 4210 8632 39120 8912
rect 4210 8232 39200 8632
rect 4210 7952 39120 8232
rect 4210 7552 39200 7952
rect 4210 7272 39120 7552
rect 4210 6872 39200 7272
rect 4210 6592 39120 6872
rect 4210 6192 39200 6592
rect 4210 5912 39120 6192
rect 4210 5512 39200 5912
rect 4210 5232 39120 5512
rect 4210 4832 39200 5232
rect 4210 4552 39120 4832
rect 4210 4152 39200 4552
rect 4210 3872 39120 4152
rect 4210 3472 39200 3872
rect 4210 3192 39120 3472
rect 4210 2792 39200 3192
rect 4210 2512 39120 2792
rect 4210 2143 39200 2512
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal3 s 39200 37272 40000 37392 6 i_clk
port 1 nsew signal input
rlabel metal3 s 39200 36592 40000 36712 6 i_rst
port 2 nsew signal input
rlabel metal2 s 37646 39200 37702 40000 6 i_wb0_cyc
port 3 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 i_wb1_cyc
port 4 nsew signal input
rlabel metal3 s 39200 35912 40000 36032 6 o_sel_sig
port 5 nsew signal output
rlabel metal3 s 39200 35232 40000 35352 6 o_wb_cyc
port 6 nsew signal output
rlabel metal3 s 39200 2592 40000 2712 6 owb_4_burst
port 7 nsew signal output
rlabel metal3 s 39200 3272 40000 3392 6 owb_8_burst
port 8 nsew signal output
rlabel metal3 s 39200 3952 40000 4072 6 owb_ack
port 9 nsew signal input
rlabel metal3 s 39200 4632 40000 4752 6 owb_adr[0]
port 10 nsew signal output
rlabel metal3 s 39200 11432 40000 11552 6 owb_adr[10]
port 11 nsew signal output
rlabel metal3 s 39200 12112 40000 12232 6 owb_adr[11]
port 12 nsew signal output
rlabel metal3 s 39200 12792 40000 12912 6 owb_adr[12]
port 13 nsew signal output
rlabel metal3 s 39200 13472 40000 13592 6 owb_adr[13]
port 14 nsew signal output
rlabel metal3 s 39200 14152 40000 14272 6 owb_adr[14]
port 15 nsew signal output
rlabel metal3 s 39200 14832 40000 14952 6 owb_adr[15]
port 16 nsew signal output
rlabel metal3 s 39200 15512 40000 15632 6 owb_adr[16]
port 17 nsew signal output
rlabel metal3 s 39200 16192 40000 16312 6 owb_adr[17]
port 18 nsew signal output
rlabel metal3 s 39200 16872 40000 16992 6 owb_adr[18]
port 19 nsew signal output
rlabel metal3 s 39200 17552 40000 17672 6 owb_adr[19]
port 20 nsew signal output
rlabel metal3 s 39200 5312 40000 5432 6 owb_adr[1]
port 21 nsew signal output
rlabel metal3 s 39200 18232 40000 18352 6 owb_adr[20]
port 22 nsew signal output
rlabel metal3 s 39200 18912 40000 19032 6 owb_adr[21]
port 23 nsew signal output
rlabel metal3 s 39200 19592 40000 19712 6 owb_adr[22]
port 24 nsew signal output
rlabel metal3 s 39200 20272 40000 20392 6 owb_adr[23]
port 25 nsew signal output
rlabel metal3 s 39200 5992 40000 6112 6 owb_adr[2]
port 26 nsew signal output
rlabel metal3 s 39200 6672 40000 6792 6 owb_adr[3]
port 27 nsew signal output
rlabel metal3 s 39200 7352 40000 7472 6 owb_adr[4]
port 28 nsew signal output
rlabel metal3 s 39200 8032 40000 8152 6 owb_adr[5]
port 29 nsew signal output
rlabel metal3 s 39200 8712 40000 8832 6 owb_adr[6]
port 30 nsew signal output
rlabel metal3 s 39200 9392 40000 9512 6 owb_adr[7]
port 31 nsew signal output
rlabel metal3 s 39200 10072 40000 10192 6 owb_adr[8]
port 32 nsew signal output
rlabel metal3 s 39200 10752 40000 10872 6 owb_adr[9]
port 33 nsew signal output
rlabel metal3 s 39200 20952 40000 21072 6 owb_err
port 34 nsew signal input
rlabel metal3 s 39200 21632 40000 21752 6 owb_o_dat[0]
port 35 nsew signal output
rlabel metal3 s 39200 28432 40000 28552 6 owb_o_dat[10]
port 36 nsew signal output
rlabel metal3 s 39200 29112 40000 29232 6 owb_o_dat[11]
port 37 nsew signal output
rlabel metal3 s 39200 29792 40000 29912 6 owb_o_dat[12]
port 38 nsew signal output
rlabel metal3 s 39200 30472 40000 30592 6 owb_o_dat[13]
port 39 nsew signal output
rlabel metal3 s 39200 31152 40000 31272 6 owb_o_dat[14]
port 40 nsew signal output
rlabel metal3 s 39200 31832 40000 31952 6 owb_o_dat[15]
port 41 nsew signal output
rlabel metal3 s 39200 22312 40000 22432 6 owb_o_dat[1]
port 42 nsew signal output
rlabel metal3 s 39200 22992 40000 23112 6 owb_o_dat[2]
port 43 nsew signal output
rlabel metal3 s 39200 23672 40000 23792 6 owb_o_dat[3]
port 44 nsew signal output
rlabel metal3 s 39200 24352 40000 24472 6 owb_o_dat[4]
port 45 nsew signal output
rlabel metal3 s 39200 25032 40000 25152 6 owb_o_dat[5]
port 46 nsew signal output
rlabel metal3 s 39200 25712 40000 25832 6 owb_o_dat[6]
port 47 nsew signal output
rlabel metal3 s 39200 26392 40000 26512 6 owb_o_dat[7]
port 48 nsew signal output
rlabel metal3 s 39200 27072 40000 27192 6 owb_o_dat[8]
port 49 nsew signal output
rlabel metal3 s 39200 27752 40000 27872 6 owb_o_dat[9]
port 50 nsew signal output
rlabel metal3 s 39200 32512 40000 32632 6 owb_sel[0]
port 51 nsew signal output
rlabel metal3 s 39200 33192 40000 33312 6 owb_sel[1]
port 52 nsew signal output
rlabel metal3 s 39200 33872 40000 33992 6 owb_stb
port 53 nsew signal output
rlabel metal3 s 39200 34552 40000 34672 6 owb_we
port 54 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 56 nsew ground bidirectional
rlabel metal2 s 2318 39200 2374 40000 6 wb0_4_burst
port 57 nsew signal input
rlabel metal2 s 3054 39200 3110 40000 6 wb0_8_burst
port 58 nsew signal input
rlabel metal2 s 3790 39200 3846 40000 6 wb0_ack
port 59 nsew signal output
rlabel metal2 s 4526 39200 4582 40000 6 wb0_adr[0]
port 60 nsew signal input
rlabel metal2 s 11886 39200 11942 40000 6 wb0_adr[10]
port 61 nsew signal input
rlabel metal2 s 12622 39200 12678 40000 6 wb0_adr[11]
port 62 nsew signal input
rlabel metal2 s 13358 39200 13414 40000 6 wb0_adr[12]
port 63 nsew signal input
rlabel metal2 s 14094 39200 14150 40000 6 wb0_adr[13]
port 64 nsew signal input
rlabel metal2 s 14830 39200 14886 40000 6 wb0_adr[14]
port 65 nsew signal input
rlabel metal2 s 15566 39200 15622 40000 6 wb0_adr[15]
port 66 nsew signal input
rlabel metal2 s 16302 39200 16358 40000 6 wb0_adr[16]
port 67 nsew signal input
rlabel metal2 s 17038 39200 17094 40000 6 wb0_adr[17]
port 68 nsew signal input
rlabel metal2 s 17774 39200 17830 40000 6 wb0_adr[18]
port 69 nsew signal input
rlabel metal2 s 18510 39200 18566 40000 6 wb0_adr[19]
port 70 nsew signal input
rlabel metal2 s 5262 39200 5318 40000 6 wb0_adr[1]
port 71 nsew signal input
rlabel metal2 s 19246 39200 19302 40000 6 wb0_adr[20]
port 72 nsew signal input
rlabel metal2 s 19982 39200 20038 40000 6 wb0_adr[21]
port 73 nsew signal input
rlabel metal2 s 20718 39200 20774 40000 6 wb0_adr[22]
port 74 nsew signal input
rlabel metal2 s 21454 39200 21510 40000 6 wb0_adr[23]
port 75 nsew signal input
rlabel metal2 s 5998 39200 6054 40000 6 wb0_adr[2]
port 76 nsew signal input
rlabel metal2 s 6734 39200 6790 40000 6 wb0_adr[3]
port 77 nsew signal input
rlabel metal2 s 7470 39200 7526 40000 6 wb0_adr[4]
port 78 nsew signal input
rlabel metal2 s 8206 39200 8262 40000 6 wb0_adr[5]
port 79 nsew signal input
rlabel metal2 s 8942 39200 8998 40000 6 wb0_adr[6]
port 80 nsew signal input
rlabel metal2 s 9678 39200 9734 40000 6 wb0_adr[7]
port 81 nsew signal input
rlabel metal2 s 10414 39200 10470 40000 6 wb0_adr[8]
port 82 nsew signal input
rlabel metal2 s 11150 39200 11206 40000 6 wb0_adr[9]
port 83 nsew signal input
rlabel metal2 s 22190 39200 22246 40000 6 wb0_err
port 84 nsew signal output
rlabel metal2 s 22926 39200 22982 40000 6 wb0_o_dat[0]
port 85 nsew signal input
rlabel metal2 s 30286 39200 30342 40000 6 wb0_o_dat[10]
port 86 nsew signal input
rlabel metal2 s 31022 39200 31078 40000 6 wb0_o_dat[11]
port 87 nsew signal input
rlabel metal2 s 31758 39200 31814 40000 6 wb0_o_dat[12]
port 88 nsew signal input
rlabel metal2 s 32494 39200 32550 40000 6 wb0_o_dat[13]
port 89 nsew signal input
rlabel metal2 s 33230 39200 33286 40000 6 wb0_o_dat[14]
port 90 nsew signal input
rlabel metal2 s 33966 39200 34022 40000 6 wb0_o_dat[15]
port 91 nsew signal input
rlabel metal2 s 23662 39200 23718 40000 6 wb0_o_dat[1]
port 92 nsew signal input
rlabel metal2 s 24398 39200 24454 40000 6 wb0_o_dat[2]
port 93 nsew signal input
rlabel metal2 s 25134 39200 25190 40000 6 wb0_o_dat[3]
port 94 nsew signal input
rlabel metal2 s 25870 39200 25926 40000 6 wb0_o_dat[4]
port 95 nsew signal input
rlabel metal2 s 26606 39200 26662 40000 6 wb0_o_dat[5]
port 96 nsew signal input
rlabel metal2 s 27342 39200 27398 40000 6 wb0_o_dat[6]
port 97 nsew signal input
rlabel metal2 s 28078 39200 28134 40000 6 wb0_o_dat[7]
port 98 nsew signal input
rlabel metal2 s 28814 39200 28870 40000 6 wb0_o_dat[8]
port 99 nsew signal input
rlabel metal2 s 29550 39200 29606 40000 6 wb0_o_dat[9]
port 100 nsew signal input
rlabel metal2 s 34702 39200 34758 40000 6 wb0_sel[0]
port 101 nsew signal input
rlabel metal2 s 35438 39200 35494 40000 6 wb0_sel[1]
port 102 nsew signal input
rlabel metal2 s 36174 39200 36230 40000 6 wb0_stb
port 103 nsew signal input
rlabel metal2 s 36910 39200 36966 40000 6 wb0_we
port 104 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wb1_4_burst
port 105 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wb1_8_burst
port 106 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wb1_ack
port 107 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 wb1_adr[0]
port 108 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wb1_adr[10]
port 109 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wb1_adr[11]
port 110 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wb1_adr[12]
port 111 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wb1_adr[13]
port 112 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wb1_adr[14]
port 113 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wb1_adr[15]
port 114 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wb1_adr[16]
port 115 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wb1_adr[17]
port 116 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wb1_adr[18]
port 117 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wb1_adr[19]
port 118 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wb1_adr[1]
port 119 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wb1_adr[20]
port 120 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wb1_adr[21]
port 121 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wb1_adr[22]
port 122 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wb1_adr[23]
port 123 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wb1_adr[2]
port 124 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wb1_adr[3]
port 125 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wb1_adr[4]
port 126 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wb1_adr[5]
port 127 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wb1_adr[6]
port 128 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wb1_adr[7]
port 129 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wb1_adr[8]
port 130 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wb1_adr[9]
port 131 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wb1_err
port 132 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 wb1_o_dat[0]
port 133 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wb1_o_dat[10]
port 134 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wb1_o_dat[11]
port 135 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wb1_o_dat[12]
port 136 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wb1_o_dat[13]
port 137 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wb1_o_dat[14]
port 138 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wb1_o_dat[15]
port 139 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wb1_o_dat[1]
port 140 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wb1_o_dat[2]
port 141 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wb1_o_dat[3]
port 142 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wb1_o_dat[4]
port 143 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wb1_o_dat[5]
port 144 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wb1_o_dat[6]
port 145 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wb1_o_dat[7]
port 146 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wb1_o_dat[8]
port 147 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wb1_o_dat[9]
port 148 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wb1_sel[0]
port 149 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wb1_sel[1]
port 150 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wb1_stb
port 151 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wb1_we
port 152 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1017362
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/wishbone_arbiter/runs/22_09_13_14_06/results/signoff/wishbone_arbiter.magic.gds
string GDS_START 104962
<< end >>

