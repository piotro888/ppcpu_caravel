magic
tech sky130B
magscale 1 2
timestamp 1663070788
<< viali >>
rect 20453 37417 20487 37451
rect 23857 37417 23891 37451
rect 30389 37417 30423 37451
rect 1777 37349 1811 37383
rect 17877 37281 17911 37315
rect 26341 37281 26375 37315
rect 34713 37281 34747 37315
rect 1593 37213 1627 37247
rect 2513 37213 2547 37247
rect 3249 37213 3283 37247
rect 4353 37213 4387 37247
rect 5089 37213 5123 37247
rect 5825 37213 5859 37247
rect 6929 37213 6963 37247
rect 7665 37213 7699 37247
rect 8401 37213 8435 37247
rect 9505 37213 9539 37247
rect 10241 37213 10275 37247
rect 10701 37213 10735 37247
rect 12081 37213 12115 37247
rect 12541 37213 12575 37247
rect 13553 37213 13587 37247
rect 14657 37213 14691 37247
rect 15393 37213 15427 37247
rect 15853 37213 15887 37247
rect 17417 37213 17451 37247
rect 18153 37213 18187 37247
rect 19625 37213 19659 37247
rect 20269 37213 20303 37247
rect 21097 37213 21131 37247
rect 22017 37213 22051 37247
rect 22661 37213 22695 37247
rect 23305 37213 23339 37247
rect 24409 37213 24443 37247
rect 25237 37213 25271 37247
rect 25881 37213 25915 37247
rect 27537 37213 27571 37247
rect 28273 37213 28307 37247
rect 29009 37213 29043 37247
rect 29837 37213 29871 37247
rect 30573 37213 30607 37247
rect 31309 37213 31343 37247
rect 32413 37213 32447 37247
rect 33149 37213 33183 37247
rect 33885 37213 33919 37247
rect 35357 37213 35391 37247
rect 37565 37213 37599 37247
rect 35624 37145 35658 37179
rect 2329 37077 2363 37111
rect 3065 37077 3099 37111
rect 4169 37077 4203 37111
rect 4905 37077 4939 37111
rect 5641 37077 5675 37111
rect 6745 37077 6779 37111
rect 7481 37077 7515 37111
rect 8217 37077 8251 37111
rect 9321 37077 9355 37111
rect 10057 37077 10091 37111
rect 10885 37077 10919 37111
rect 11897 37077 11931 37111
rect 12725 37077 12759 37111
rect 13369 37077 13403 37111
rect 14473 37077 14507 37111
rect 15209 37077 15243 37111
rect 16037 37077 16071 37111
rect 17233 37077 17267 37111
rect 19809 37077 19843 37111
rect 20913 37077 20947 37111
rect 21833 37077 21867 37111
rect 22477 37077 22511 37111
rect 23121 37077 23155 37111
rect 24593 37077 24627 37111
rect 25053 37077 25087 37111
rect 25697 37077 25731 37111
rect 27353 37077 27387 37111
rect 28089 37077 28123 37111
rect 28825 37077 28859 37111
rect 29653 37077 29687 37111
rect 31125 37077 31159 37111
rect 32229 37077 32263 37111
rect 32965 37077 32999 37111
rect 33701 37077 33735 37111
rect 36737 37077 36771 37111
rect 37381 37077 37415 37111
rect 38117 37077 38151 37111
rect 1869 36873 1903 36907
rect 2513 36873 2547 36907
rect 4721 36873 4755 36907
rect 6469 36873 6503 36907
rect 8033 36873 8067 36907
rect 9137 36873 9171 36907
rect 10793 36873 10827 36907
rect 12449 36873 12483 36907
rect 14105 36873 14139 36907
rect 15761 36873 15795 36907
rect 16865 36873 16899 36907
rect 19993 36873 20027 36907
rect 20821 36873 20855 36907
rect 20913 36873 20947 36907
rect 21281 36873 21315 36907
rect 23673 36873 23707 36907
rect 24133 36873 24167 36907
rect 30757 36873 30791 36907
rect 35909 36873 35943 36907
rect 37381 36873 37415 36907
rect 3065 36805 3099 36839
rect 3617 36805 3651 36839
rect 13553 36805 13587 36839
rect 19257 36805 19291 36839
rect 29938 36805 29972 36839
rect 33250 36805 33284 36839
rect 35090 36805 35124 36839
rect 4905 36737 4939 36771
rect 6653 36737 6687 36771
rect 8217 36737 8251 36771
rect 9321 36737 9355 36771
rect 10977 36737 11011 36771
rect 12633 36737 12667 36771
rect 14289 36737 14323 36771
rect 15209 36737 15243 36771
rect 15945 36737 15979 36771
rect 17049 36737 17083 36771
rect 17509 36737 17543 36771
rect 18153 36737 18187 36771
rect 19165 36737 19199 36771
rect 21833 36737 21867 36771
rect 23305 36737 23339 36771
rect 25246 36737 25280 36771
rect 26157 36737 26191 36771
rect 28098 36737 28132 36771
rect 30941 36737 30975 36771
rect 36093 36737 36127 36771
rect 37565 36737 37599 36771
rect 19441 36669 19475 36703
rect 20729 36669 20763 36703
rect 23029 36669 23063 36703
rect 23213 36669 23247 36703
rect 25513 36669 25547 36703
rect 28365 36669 28399 36703
rect 30205 36669 30239 36703
rect 33517 36669 33551 36703
rect 35357 36669 35391 36703
rect 3801 36601 3835 36635
rect 18797 36601 18831 36635
rect 22017 36601 22051 36635
rect 28825 36601 28859 36635
rect 32137 36601 32171 36635
rect 5825 36533 5859 36567
rect 7389 36533 7423 36567
rect 10241 36533 10275 36567
rect 11897 36533 11931 36567
rect 17693 36533 17727 36567
rect 18337 36533 18371 36567
rect 25973 36533 26007 36567
rect 26985 36533 27019 36567
rect 31401 36533 31435 36567
rect 33977 36533 34011 36567
rect 36645 36533 36679 36567
rect 14473 36329 14507 36363
rect 16957 36329 16991 36363
rect 19441 36329 19475 36363
rect 20177 36329 20211 36363
rect 22753 36329 22787 36363
rect 29561 36329 29595 36363
rect 37197 36329 37231 36363
rect 6837 36261 6871 36295
rect 16405 36261 16439 36295
rect 18705 36261 18739 36295
rect 22109 36261 22143 36295
rect 23397 36261 23431 36295
rect 37933 36261 37967 36295
rect 2697 36193 2731 36227
rect 9505 36193 9539 36227
rect 15301 36193 15335 36227
rect 20729 36193 20763 36227
rect 21557 36193 21591 36227
rect 21649 36193 21683 36227
rect 33793 36193 33827 36227
rect 7389 36125 7423 36159
rect 10425 36125 10459 36159
rect 13553 36125 13587 36159
rect 17509 36125 17543 36159
rect 18521 36125 18555 36159
rect 19349 36125 19383 36159
rect 22569 36125 22603 36159
rect 23213 36125 23247 36159
rect 24409 36125 24443 36159
rect 26525 36125 26559 36159
rect 28558 36125 28592 36159
rect 28825 36125 28859 36159
rect 30205 36125 30239 36159
rect 35173 36125 35207 36159
rect 37013 36125 37047 36159
rect 37749 36125 37783 36159
rect 5641 36057 5675 36091
rect 11161 36057 11195 36091
rect 18061 36057 18095 36091
rect 20637 36057 20671 36091
rect 21741 36057 21775 36091
rect 26258 36057 26292 36091
rect 30450 36057 30484 36091
rect 33526 36057 33560 36091
rect 35440 36057 35474 36091
rect 4537 35989 4571 36023
rect 5089 35989 5123 36023
rect 8401 35989 8435 36023
rect 12173 35989 12207 36023
rect 12817 35989 12851 36023
rect 15853 35989 15887 36023
rect 20545 35989 20579 36023
rect 24593 35989 24627 36023
rect 25145 35989 25179 36023
rect 27445 35989 27479 36023
rect 31585 35989 31619 36023
rect 32413 35989 32447 36023
rect 36553 35989 36587 36023
rect 17233 35785 17267 35819
rect 17877 35785 17911 35819
rect 18521 35785 18555 35819
rect 21097 35785 21131 35819
rect 22109 35785 22143 35819
rect 22569 35785 22603 35819
rect 23765 35785 23799 35819
rect 26985 35785 27019 35819
rect 30573 35785 30607 35819
rect 32873 35785 32907 35819
rect 33609 35785 33643 35819
rect 34345 35785 34379 35819
rect 36185 35785 36219 35819
rect 37841 35785 37875 35819
rect 13369 35717 13403 35751
rect 19257 35717 19291 35751
rect 23305 35717 23339 35751
rect 13737 35649 13771 35683
rect 13829 35649 13863 35683
rect 14565 35649 14599 35683
rect 15209 35649 15243 35683
rect 19349 35649 19383 35683
rect 20177 35649 20211 35683
rect 22201 35649 22235 35683
rect 23397 35649 23431 35683
rect 25338 35649 25372 35683
rect 25605 35649 25639 35683
rect 26249 35649 26283 35683
rect 27169 35649 27203 35683
rect 29294 35649 29328 35683
rect 33057 35649 33091 35683
rect 33793 35649 33827 35683
rect 34529 35649 34563 35683
rect 36369 35649 36403 35683
rect 38025 35649 38059 35683
rect 13461 35581 13495 35615
rect 14749 35581 14783 35615
rect 14841 35581 14875 35615
rect 19165 35581 19199 35615
rect 21925 35581 21959 35615
rect 23121 35581 23155 35615
rect 27629 35581 27663 35615
rect 29561 35581 29595 35615
rect 24225 35513 24259 35547
rect 8585 35445 8619 35479
rect 9689 35445 9723 35479
rect 13553 35445 13587 35479
rect 19717 35445 19751 35479
rect 20361 35445 20395 35479
rect 26065 35445 26099 35479
rect 28181 35445 28215 35479
rect 30113 35445 30147 35479
rect 31125 35445 31159 35479
rect 32137 35445 32171 35479
rect 34989 35445 35023 35479
rect 35633 35445 35667 35479
rect 15393 35241 15427 35275
rect 19349 35241 19383 35275
rect 26709 35241 26743 35275
rect 27905 35241 27939 35275
rect 14473 35173 14507 35207
rect 22753 35173 22787 35207
rect 25881 35173 25915 35207
rect 31401 35173 31435 35207
rect 16405 35105 16439 35139
rect 17233 35105 17267 35139
rect 14749 35037 14783 35071
rect 15393 35037 15427 35071
rect 15577 35037 15611 35071
rect 16221 35037 16255 35071
rect 16313 35037 16347 35071
rect 16497 35037 16531 35071
rect 16681 35037 16715 35071
rect 19809 35037 19843 35071
rect 21005 35037 21039 35071
rect 23213 35037 23247 35071
rect 23857 35037 23891 35071
rect 24685 35037 24719 35071
rect 25329 35037 25363 35071
rect 26893 35037 26927 35071
rect 27353 35037 27387 35071
rect 30021 35037 30055 35071
rect 33517 35037 33551 35071
rect 34069 35037 34103 35071
rect 36093 35037 36127 35071
rect 36737 35037 36771 35071
rect 14473 34969 14507 35003
rect 30266 34969 30300 35003
rect 33250 34969 33284 35003
rect 35826 34969 35860 35003
rect 37004 34969 37038 35003
rect 12357 34901 12391 34935
rect 14657 34901 14691 34935
rect 16037 34901 16071 34935
rect 19993 34901 20027 34935
rect 21097 34901 21131 34935
rect 21833 34901 21867 34935
rect 24501 34901 24535 34935
rect 25145 34901 25179 34935
rect 28457 34901 28491 34935
rect 32137 34901 32171 34935
rect 34713 34901 34747 34935
rect 38117 34901 38151 34935
rect 9597 34697 9631 34731
rect 10885 34697 10919 34731
rect 12087 34697 12121 34731
rect 14565 34697 14599 34731
rect 21005 34697 21039 34731
rect 22017 34697 22051 34731
rect 22753 34697 22787 34731
rect 23397 34697 23431 34731
rect 24317 34697 24351 34731
rect 26249 34697 26283 34731
rect 26985 34697 27019 34731
rect 29101 34697 29135 34731
rect 10057 34629 10091 34663
rect 14749 34629 14783 34663
rect 15669 34629 15703 34663
rect 34170 34629 34204 34663
rect 10241 34561 10275 34595
rect 10333 34561 10367 34595
rect 11989 34561 12023 34595
rect 12173 34561 12207 34595
rect 12265 34561 12299 34595
rect 12909 34561 12943 34595
rect 13093 34561 13127 34595
rect 13553 34561 13587 34595
rect 14933 34561 14967 34595
rect 20637 34561 20671 34595
rect 21833 34561 21867 34595
rect 22569 34561 22603 34595
rect 23213 34561 23247 34595
rect 25430 34561 25464 34595
rect 25697 34561 25731 34595
rect 28098 34561 28132 34595
rect 28365 34561 28399 34595
rect 30214 34561 30248 34595
rect 30481 34561 30515 34595
rect 13645 34493 13679 34527
rect 19625 34493 19659 34527
rect 20453 34493 20487 34527
rect 20545 34493 20579 34527
rect 34437 34493 34471 34527
rect 35909 34493 35943 34527
rect 37289 34493 37323 34527
rect 10057 34425 10091 34459
rect 36277 34425 36311 34459
rect 37841 34425 37875 34459
rect 13001 34357 13035 34391
rect 33057 34357 33091 34391
rect 36369 34357 36403 34391
rect 10609 34153 10643 34187
rect 15209 34153 15243 34187
rect 16681 34153 16715 34187
rect 22201 34153 22235 34187
rect 22937 34153 22971 34187
rect 24961 34153 24995 34187
rect 25605 34153 25639 34187
rect 29009 34153 29043 34187
rect 36093 34153 36127 34187
rect 12265 34085 12299 34119
rect 12817 34085 12851 34119
rect 26709 34085 26743 34119
rect 10057 34017 10091 34051
rect 11713 34017 11747 34051
rect 11989 34017 12023 34051
rect 20913 34017 20947 34051
rect 23489 34017 23523 34051
rect 24501 34017 24535 34051
rect 26065 34017 26099 34051
rect 28089 34017 28123 34051
rect 9229 33949 9263 33983
rect 9413 33949 9447 33983
rect 11529 33949 11563 33983
rect 12265 33949 12299 33983
rect 13185 33949 13219 33983
rect 14105 33949 14139 33983
rect 17693 33949 17727 33983
rect 17856 33949 17890 33983
rect 17956 33943 17990 33977
rect 18061 33949 18095 33983
rect 21373 33949 21407 33983
rect 22017 33949 22051 33983
rect 23397 33949 23431 33983
rect 27822 33949 27856 33983
rect 34713 33949 34747 33983
rect 36737 33949 36771 33983
rect 13001 33881 13035 33915
rect 15025 33881 15059 33915
rect 15225 33881 15259 33915
rect 16405 33881 16439 33915
rect 16589 33881 16623 33915
rect 18337 33881 18371 33915
rect 19349 33881 19383 33915
rect 32965 33881 32999 33915
rect 34958 33881 34992 33915
rect 37004 33881 37038 33915
rect 9413 33813 9447 33847
rect 10149 33813 10183 33847
rect 10241 33813 10275 33847
rect 14289 33813 14323 33847
rect 15393 33813 15427 33847
rect 21557 33813 21591 33847
rect 23305 33813 23339 33847
rect 31677 33813 31711 33847
rect 38117 33813 38151 33847
rect 8769 33609 8803 33643
rect 10793 33609 10827 33643
rect 13001 33609 13035 33643
rect 19993 33609 20027 33643
rect 20453 33609 20487 33643
rect 21833 33609 21867 33643
rect 23029 33609 23063 33643
rect 23489 33609 23523 33643
rect 36277 33609 36311 33643
rect 9413 33541 9447 33575
rect 22293 33541 22327 33575
rect 9321 33473 9355 33507
rect 9505 33473 9539 33507
rect 10425 33473 10459 33507
rect 10609 33473 10643 33507
rect 11529 33473 11563 33507
rect 12725 33473 12759 33507
rect 12817 33473 12851 33507
rect 13921 33473 13955 33507
rect 16681 33473 16715 33507
rect 18245 33473 18279 33507
rect 20085 33473 20119 33507
rect 20913 33473 20947 33507
rect 22201 33473 22235 33507
rect 23397 33473 23431 33507
rect 24317 33473 24351 33507
rect 28641 33473 28675 33507
rect 33793 33473 33827 33507
rect 36093 33473 36127 33507
rect 19901 33405 19935 33439
rect 22477 33405 22511 33439
rect 23581 33405 23615 33439
rect 35541 33405 35575 33439
rect 16865 33337 16899 33371
rect 10517 33269 10551 33303
rect 14105 33269 14139 33303
rect 14841 33269 14875 33303
rect 17601 33269 17635 33303
rect 18429 33269 18463 33303
rect 29929 33269 29963 33303
rect 9781 33065 9815 33099
rect 12725 33065 12759 33099
rect 18429 33065 18463 33099
rect 28273 33065 28307 33099
rect 22753 32997 22787 33031
rect 23305 32997 23339 33031
rect 24409 32997 24443 33031
rect 30481 32997 30515 33031
rect 17785 32929 17819 32963
rect 17969 32929 18003 32963
rect 12817 32861 12851 32895
rect 25789 32861 25823 32895
rect 26893 32861 26927 32895
rect 31594 32861 31628 32895
rect 31861 32861 31895 32895
rect 33701 32861 33735 32895
rect 13277 32793 13311 32827
rect 18061 32793 18095 32827
rect 19349 32793 19383 32827
rect 25522 32793 25556 32827
rect 27138 32793 27172 32827
rect 33434 32793 33468 32827
rect 14197 32725 14231 32759
rect 32321 32725 32355 32759
rect 12449 32521 12483 32555
rect 36369 32521 36403 32555
rect 13185 32453 13219 32487
rect 14013 32453 14047 32487
rect 25798 32453 25832 32487
rect 12265 32385 12299 32419
rect 13461 32385 13495 32419
rect 13921 32385 13955 32419
rect 14381 32385 14415 32419
rect 18245 32385 18279 32419
rect 18981 32385 19015 32419
rect 19165 32385 19199 32419
rect 19717 32385 19751 32419
rect 22661 32385 22695 32419
rect 26065 32385 26099 32419
rect 28926 32385 28960 32419
rect 29909 32385 29943 32419
rect 35245 32385 35279 32419
rect 13185 32317 13219 32351
rect 14289 32317 14323 32351
rect 14933 32317 14967 32351
rect 18797 32317 18831 32351
rect 29193 32317 29227 32351
rect 29653 32317 29687 32351
rect 34989 32317 35023 32351
rect 19901 32249 19935 32283
rect 22845 32249 22879 32283
rect 31033 32249 31067 32283
rect 13369 32181 13403 32215
rect 14197 32181 14231 32215
rect 21833 32181 21867 32215
rect 24685 32181 24719 32215
rect 27813 32181 27847 32215
rect 13553 31977 13587 32011
rect 14565 31977 14599 32011
rect 16865 31977 16899 32011
rect 22201 31977 22235 32011
rect 29653 31977 29687 32011
rect 34805 31977 34839 32011
rect 38117 31977 38151 32011
rect 21557 31909 21591 31943
rect 24409 31909 24443 31943
rect 31309 31909 31343 31943
rect 15945 31841 15979 31875
rect 16221 31841 16255 31875
rect 20913 31841 20947 31875
rect 21097 31841 21131 31875
rect 25789 31841 25823 31875
rect 36737 31841 36771 31875
rect 15853 31773 15887 31807
rect 16681 31773 16715 31807
rect 19349 31773 19383 31807
rect 22017 31773 22051 31807
rect 22937 31773 22971 31807
rect 25522 31773 25556 31807
rect 32689 31773 32723 31807
rect 36993 31773 37027 31807
rect 21189 31705 21223 31739
rect 32422 31705 32456 31739
rect 23121 31637 23155 31671
rect 30757 31637 30791 31671
rect 35265 31637 35299 31671
rect 22109 31365 22143 31399
rect 25430 31365 25464 31399
rect 27230 31365 27264 31399
rect 34253 31365 34287 31399
rect 16681 31297 16715 31331
rect 18705 31297 18739 31331
rect 20453 31297 20487 31331
rect 22201 31297 22235 31331
rect 23029 31297 23063 31331
rect 25697 31297 25731 31331
rect 26985 31297 27019 31331
rect 30214 31297 30248 31331
rect 30481 31297 30515 31331
rect 34713 31297 34747 31331
rect 34969 31297 35003 31331
rect 18613 31229 18647 31263
rect 19073 31229 19107 31263
rect 21925 31229 21959 31263
rect 16865 31161 16899 31195
rect 17969 31093 18003 31127
rect 20637 31093 20671 31127
rect 22569 31093 22603 31127
rect 24317 31093 24351 31127
rect 28365 31093 28399 31127
rect 29101 31093 29135 31127
rect 32965 31093 32999 31127
rect 36093 31093 36127 31127
rect 12173 30889 12207 30923
rect 18429 30889 18463 30923
rect 20913 30889 20947 30923
rect 30941 30889 30975 30923
rect 36461 30889 36495 30923
rect 17049 30753 17083 30787
rect 17141 30753 17175 30787
rect 26065 30753 26099 30787
rect 11805 30685 11839 30719
rect 11989 30685 12023 30719
rect 12633 30685 12667 30719
rect 18153 30685 18187 30719
rect 18245 30685 18279 30719
rect 20085 30685 20119 30719
rect 20545 30685 20579 30719
rect 20729 30685 20763 30719
rect 27813 30685 27847 30719
rect 32321 30685 32355 30719
rect 35081 30685 35115 30719
rect 17233 30617 17267 30651
rect 32054 30617 32088 30651
rect 35348 30617 35382 30651
rect 12817 30549 12851 30583
rect 17601 30549 17635 30583
rect 11897 30277 11931 30311
rect 15485 30277 15519 30311
rect 22385 30277 22419 30311
rect 25522 30277 25556 30311
rect 11713 30209 11747 30243
rect 13737 30209 13771 30243
rect 14381 30209 14415 30243
rect 15301 30209 15335 30243
rect 17509 30209 17543 30243
rect 28190 30209 28224 30243
rect 29173 30209 29207 30243
rect 34630 30209 34664 30243
rect 11529 30141 11563 30175
rect 15117 30141 15151 30175
rect 25789 30141 25823 30175
rect 28457 30141 28491 30175
rect 28917 30141 28951 30175
rect 34897 30141 34931 30175
rect 17693 30073 17727 30107
rect 13093 30005 13127 30039
rect 14289 30005 14323 30039
rect 18245 30005 18279 30039
rect 21925 30005 21959 30039
rect 24409 30005 24443 30039
rect 27077 30005 27111 30039
rect 30297 30005 30331 30039
rect 33517 30005 33551 30039
rect 12265 29801 12299 29835
rect 16497 29801 16531 29835
rect 36277 29801 36311 29835
rect 38117 29801 38151 29835
rect 13553 29733 13587 29767
rect 22017 29733 22051 29767
rect 12817 29665 12851 29699
rect 15761 29665 15795 29699
rect 21300 29665 21334 29699
rect 21833 29665 21867 29699
rect 32045 29665 32079 29699
rect 12725 29597 12759 29631
rect 14105 29597 14139 29631
rect 15577 29597 15611 29631
rect 17049 29597 17083 29631
rect 21097 29597 21131 29631
rect 22108 29597 22142 29631
rect 22569 29597 22603 29631
rect 23305 29597 23339 29631
rect 25789 29597 25823 29631
rect 34897 29597 34931 29631
rect 36737 29597 36771 29631
rect 21373 29529 21407 29563
rect 21833 29529 21867 29563
rect 25522 29529 25556 29563
rect 31778 29529 31812 29563
rect 35164 29529 35198 29563
rect 36982 29529 37016 29563
rect 12633 29461 12667 29495
rect 14289 29461 14323 29495
rect 15209 29461 15243 29495
rect 15669 29461 15703 29495
rect 17233 29461 17267 29495
rect 21189 29461 21223 29495
rect 22753 29461 22787 29495
rect 24409 29461 24443 29495
rect 30665 29461 30699 29495
rect 10241 29257 10275 29291
rect 13185 29257 13219 29291
rect 15577 29257 15611 29291
rect 20821 29189 20855 29223
rect 20913 29189 20947 29223
rect 25522 29189 25556 29223
rect 12173 29121 12207 29155
rect 13001 29121 13035 29155
rect 15393 29121 15427 29155
rect 19533 29121 19567 29155
rect 21833 29121 21867 29155
rect 22017 29121 22051 29155
rect 22201 29121 22235 29155
rect 29110 29121 29144 29155
rect 29377 29121 29411 29155
rect 33986 29121 34020 29155
rect 34253 29121 34287 29155
rect 15209 29053 15243 29087
rect 20729 29053 20763 29087
rect 22661 29053 22695 29087
rect 25789 29053 25823 29087
rect 10793 28985 10827 29019
rect 12357 28985 12391 29019
rect 16037 28985 16071 29019
rect 19717 28985 19751 29019
rect 24409 28985 24443 29019
rect 27997 28985 28031 29019
rect 32873 28985 32907 29019
rect 9689 28917 9723 28951
rect 11529 28917 11563 28951
rect 21281 28917 21315 28951
rect 14105 28713 14139 28747
rect 17417 28713 17451 28747
rect 27629 28713 27663 28747
rect 30941 28713 30975 28747
rect 38117 28713 38151 28747
rect 25053 28645 25087 28679
rect 9689 28577 9723 28611
rect 10793 28577 10827 28611
rect 15761 28577 15795 28611
rect 21833 28577 21867 28611
rect 29009 28577 29043 28611
rect 32321 28577 32355 28611
rect 9505 28509 9539 28543
rect 10701 28509 10735 28543
rect 11621 28509 11655 28543
rect 14289 28509 14323 28543
rect 14473 28509 14507 28543
rect 17049 28509 17083 28543
rect 17233 28509 17267 28543
rect 21189 28509 21223 28543
rect 26433 28509 26467 28543
rect 36737 28509 36771 28543
rect 10609 28441 10643 28475
rect 12357 28441 12391 28475
rect 15025 28441 15059 28475
rect 15209 28441 15243 28475
rect 26166 28441 26200 28475
rect 28742 28441 28776 28475
rect 32054 28441 32088 28475
rect 36982 28441 37016 28475
rect 9045 28373 9079 28407
rect 9413 28373 9447 28407
rect 10241 28373 10275 28407
rect 11805 28373 11839 28407
rect 12909 28373 12943 28407
rect 16221 28373 16255 28407
rect 21373 28373 21407 28407
rect 9965 28169 9999 28203
rect 12265 28169 12299 28203
rect 12725 28169 12759 28203
rect 15393 28169 15427 28203
rect 15761 28169 15795 28203
rect 19165 28169 19199 28203
rect 25154 28101 25188 28135
rect 35182 28101 35216 28135
rect 9045 28033 9079 28067
rect 9229 28033 9263 28067
rect 9781 28033 9815 28067
rect 10609 28033 10643 28067
rect 11897 28033 11931 28067
rect 12081 28033 12115 28067
rect 12909 28033 12943 28067
rect 15853 28033 15887 28067
rect 16681 28033 16715 28067
rect 18981 28033 19015 28067
rect 29754 28033 29788 28067
rect 30021 28033 30055 28067
rect 8861 27965 8895 27999
rect 10425 27965 10459 27999
rect 13093 27965 13127 27999
rect 15945 27965 15979 27999
rect 18797 27965 18831 27999
rect 25421 27965 25455 27999
rect 35449 27965 35483 27999
rect 16865 27897 16899 27931
rect 24041 27897 24075 27931
rect 10793 27829 10827 27863
rect 13553 27829 13587 27863
rect 14933 27829 14967 27863
rect 20269 27829 20303 27863
rect 28641 27829 28675 27863
rect 34069 27829 34103 27863
rect 11253 27625 11287 27659
rect 11989 27625 12023 27659
rect 15669 27557 15703 27591
rect 18061 27557 18095 27591
rect 18705 27557 18739 27591
rect 19257 27557 19291 27591
rect 32781 27557 32815 27591
rect 35633 27557 35667 27591
rect 10885 27489 10919 27523
rect 12633 27489 12667 27523
rect 14289 27489 14323 27523
rect 15301 27489 15335 27523
rect 20729 27489 20763 27523
rect 27721 27489 27755 27523
rect 11069 27421 11103 27455
rect 12357 27421 12391 27455
rect 13277 27421 13311 27455
rect 15485 27421 15519 27455
rect 16405 27421 16439 27455
rect 17877 27421 17911 27455
rect 18521 27421 18555 27455
rect 20361 27421 20395 27455
rect 20545 27421 20579 27455
rect 21649 27421 21683 27455
rect 22293 27421 22327 27455
rect 25789 27421 25823 27455
rect 34161 27421 34195 27455
rect 37013 27421 37047 27455
rect 12449 27353 12483 27387
rect 14381 27353 14415 27387
rect 25522 27353 25556 27387
rect 27454 27353 27488 27387
rect 33894 27353 33928 27387
rect 36746 27353 36780 27387
rect 14473 27285 14507 27319
rect 14841 27285 14875 27319
rect 19901 27285 19935 27319
rect 21833 27285 21867 27319
rect 22477 27285 22511 27319
rect 24409 27285 24443 27319
rect 26341 27285 26375 27319
rect 12357 27081 12391 27115
rect 12725 27081 12759 27115
rect 13553 27081 13587 27115
rect 17785 27081 17819 27115
rect 20821 27081 20855 27115
rect 32137 27081 32171 27115
rect 35357 27081 35391 27115
rect 15301 27013 15335 27047
rect 29990 27013 30024 27047
rect 8585 26945 8619 26979
rect 9413 26945 9447 26979
rect 9597 26945 9631 26979
rect 10057 26945 10091 26979
rect 11621 26945 11655 26979
rect 12817 26945 12851 26979
rect 14381 26945 14415 26979
rect 14565 26945 14599 26979
rect 17601 26945 17635 26979
rect 18889 26945 18923 26979
rect 19073 26945 19107 26979
rect 19257 26945 19291 26979
rect 19717 26945 19751 26979
rect 20545 26945 20579 26979
rect 20637 26945 20671 26979
rect 22109 26945 22143 26979
rect 25522 26945 25556 26979
rect 28098 26945 28132 26979
rect 28365 26945 28399 26979
rect 29745 26945 29779 26979
rect 33250 26945 33284 26979
rect 33517 26945 33551 26979
rect 33977 26945 34011 26979
rect 34233 26945 34267 26979
rect 8401 26877 8435 26911
rect 9229 26877 9263 26911
rect 12909 26877 12943 26911
rect 17417 26877 17451 26911
rect 21925 26877 21959 26911
rect 25789 26877 25823 26911
rect 10241 26809 10275 26843
rect 11805 26809 11839 26843
rect 26985 26809 27019 26843
rect 8769 26741 8803 26775
rect 14749 26741 14783 26775
rect 15945 26741 15979 26775
rect 16957 26741 16991 26775
rect 18337 26741 18371 26775
rect 19901 26741 19935 26775
rect 22293 26741 22327 26775
rect 22845 26741 22879 26775
rect 24409 26741 24443 26775
rect 31125 26741 31159 26775
rect 9137 26537 9171 26571
rect 11253 26537 11287 26571
rect 17141 26537 17175 26571
rect 20453 26537 20487 26571
rect 21189 26537 21223 26571
rect 37657 26537 37691 26571
rect 11897 26469 11931 26503
rect 14933 26469 14967 26503
rect 18613 26469 18647 26503
rect 9689 26401 9723 26435
rect 10885 26401 10919 26435
rect 17969 26401 18003 26435
rect 19441 26401 19475 26435
rect 21741 26401 21775 26435
rect 32965 26401 32999 26435
rect 9505 26333 9539 26367
rect 10333 26333 10367 26367
rect 11069 26333 11103 26367
rect 11713 26333 11747 26367
rect 14749 26333 14783 26367
rect 16773 26333 16807 26367
rect 16957 26333 16991 26367
rect 18245 26333 18279 26367
rect 21557 26333 21591 26367
rect 27813 26333 27847 26367
rect 31217 26333 31251 26367
rect 35357 26333 35391 26367
rect 9597 26265 9631 26299
rect 13185 26265 13219 26299
rect 16313 26265 16347 26299
rect 18153 26265 18187 26299
rect 19533 26265 19567 26299
rect 21649 26265 21683 26299
rect 22385 26265 22419 26299
rect 23029 26265 23063 26299
rect 26249 26265 26283 26299
rect 36369 26265 36403 26299
rect 19625 26197 19659 26231
rect 19993 26197 20027 26231
rect 35541 26197 35575 26231
rect 9321 25993 9355 26027
rect 16037 25993 16071 26027
rect 16681 25993 16715 26027
rect 18337 25993 18371 26027
rect 29101 25993 29135 26027
rect 32137 25993 32171 26027
rect 36737 25993 36771 26027
rect 37841 25993 37875 26027
rect 17049 25925 17083 25959
rect 30389 25925 30423 25959
rect 35624 25925 35658 25959
rect 9137 25857 9171 25891
rect 20729 25857 20763 25891
rect 22201 25857 22235 25891
rect 25246 25857 25280 25891
rect 33261 25857 33295 25891
rect 33517 25857 33551 25891
rect 38025 25857 38059 25891
rect 17141 25789 17175 25823
rect 17233 25789 17267 25823
rect 21833 25789 21867 25823
rect 22293 25789 22327 25823
rect 25513 25789 25547 25823
rect 35357 25789 35391 25823
rect 19901 25721 19935 25755
rect 24133 25721 24167 25755
rect 10149 25653 10183 25687
rect 10793 25653 10827 25687
rect 12449 25653 12483 25687
rect 15577 25653 15611 25687
rect 18889 25653 18923 25687
rect 20453 25653 20487 25687
rect 8953 25449 8987 25483
rect 11621 25449 11655 25483
rect 12909 25449 12943 25483
rect 15853 25449 15887 25483
rect 18705 25449 18739 25483
rect 26249 25449 26283 25483
rect 33885 25449 33919 25483
rect 35357 25449 35391 25483
rect 10241 25381 10275 25415
rect 13461 25381 13495 25415
rect 22661 25381 22695 25415
rect 24409 25381 24443 25415
rect 34897 25381 34931 25415
rect 9597 25313 9631 25347
rect 12265 25313 12299 25347
rect 15209 25313 15243 25347
rect 17141 25313 17175 25347
rect 18061 25313 18095 25347
rect 29561 25313 29595 25347
rect 36737 25313 36771 25347
rect 9321 25245 9355 25279
rect 11989 25245 12023 25279
rect 15485 25245 15519 25279
rect 17417 25245 17451 25279
rect 18337 25245 18371 25279
rect 22477 25245 22511 25279
rect 25522 25245 25556 25279
rect 25789 25245 25823 25279
rect 27629 25245 27663 25279
rect 29817 25245 29851 25279
rect 32781 25245 32815 25279
rect 33701 25245 33735 25279
rect 34713 25245 34747 25279
rect 35541 25245 35575 25279
rect 35725 25245 35759 25279
rect 36185 25245 36219 25279
rect 9413 25177 9447 25211
rect 15393 25177 15427 25211
rect 16589 25177 16623 25211
rect 19533 25177 19567 25211
rect 23213 25177 23247 25211
rect 27362 25177 27396 25211
rect 32514 25177 32548 25211
rect 36982 25177 37016 25211
rect 10701 25109 10735 25143
rect 12081 25109 12115 25143
rect 14105 25109 14139 25143
rect 18245 25109 18279 25143
rect 19993 25109 20027 25143
rect 20637 25109 20671 25143
rect 21097 25109 21131 25143
rect 21833 25109 21867 25143
rect 23765 25109 23799 25143
rect 30941 25109 30975 25143
rect 31401 25109 31435 25143
rect 38117 25109 38151 25143
rect 9873 24905 9907 24939
rect 13645 24905 13679 24939
rect 14841 24905 14875 24939
rect 15669 24905 15703 24939
rect 20453 24905 20487 24939
rect 37749 24905 37783 24939
rect 11897 24837 11931 24871
rect 17601 24837 17635 24871
rect 14933 24769 14967 24803
rect 16681 24769 16715 24803
rect 19073 24769 19107 24803
rect 22201 24769 22235 24803
rect 22385 24769 22419 24803
rect 22569 24769 22603 24803
rect 23121 24769 23155 24803
rect 28834 24769 28868 24803
rect 29101 24769 29135 24803
rect 29561 24769 29595 24803
rect 31217 24769 31251 24803
rect 33057 24769 33091 24803
rect 35173 24769 35207 24803
rect 36001 24769 36035 24803
rect 37657 24769 37691 24803
rect 11989 24701 12023 24735
rect 12173 24701 12207 24735
rect 13737 24701 13771 24735
rect 13829 24701 13863 24735
rect 15025 24701 15059 24735
rect 17693 24701 17727 24735
rect 17877 24701 17911 24735
rect 18521 24701 18555 24735
rect 19257 24701 19291 24735
rect 20177 24701 20211 24735
rect 20361 24701 20395 24735
rect 24317 24701 24351 24735
rect 37473 24701 37507 24735
rect 11529 24633 11563 24667
rect 13277 24633 13311 24667
rect 14473 24633 14507 24667
rect 17233 24633 17267 24667
rect 20821 24633 20855 24667
rect 27721 24633 27755 24667
rect 29745 24633 29779 24667
rect 31401 24633 31435 24667
rect 33241 24633 33275 24667
rect 35357 24633 35391 24667
rect 36185 24633 36219 24667
rect 12817 24565 12851 24599
rect 23305 24565 23339 24599
rect 23765 24565 23799 24599
rect 30205 24565 30239 24599
rect 32137 24565 32171 24599
rect 33701 24565 33735 24599
rect 34345 24565 34379 24599
rect 36737 24565 36771 24599
rect 38117 24565 38151 24599
rect 14289 24361 14323 24395
rect 17785 24361 17819 24395
rect 21189 24361 21223 24395
rect 22109 24361 22143 24395
rect 28089 24361 28123 24395
rect 29561 24361 29595 24395
rect 32137 24361 32171 24395
rect 35541 24361 35575 24395
rect 36553 24361 36587 24395
rect 38117 24361 38151 24395
rect 20453 24293 20487 24327
rect 25053 24293 25087 24327
rect 28825 24293 28859 24327
rect 30573 24293 30607 24327
rect 37013 24293 37047 24327
rect 18337 24225 18371 24259
rect 19625 24225 19659 24259
rect 22753 24225 22787 24259
rect 33425 24225 33459 24259
rect 18521 24157 18555 24191
rect 19809 24157 19843 24191
rect 19993 24157 20027 24191
rect 21005 24157 21039 24191
rect 27905 24157 27939 24191
rect 28641 24157 28675 24191
rect 29745 24157 29779 24191
rect 29837 24157 29871 24191
rect 30389 24157 30423 24191
rect 31033 24157 31067 24191
rect 31769 24157 31803 24191
rect 31953 24157 31987 24191
rect 33149 24157 33183 24191
rect 34713 24157 34747 24191
rect 34897 24157 34931 24191
rect 35725 24157 35759 24191
rect 36369 24157 36403 24191
rect 37749 24157 37783 24191
rect 37933 24157 37967 24191
rect 22569 24089 22603 24123
rect 35081 24089 35115 24123
rect 12541 24021 12575 24055
rect 15301 24021 15335 24055
rect 17325 24021 17359 24055
rect 18705 24021 18739 24055
rect 22477 24021 22511 24055
rect 23397 24021 23431 24055
rect 24501 24021 24535 24055
rect 25605 24021 25639 24055
rect 31217 24021 31251 24055
rect 32781 24021 32815 24055
rect 33241 24021 33275 24055
rect 34069 24021 34103 24055
rect 17417 23817 17451 23851
rect 18889 23817 18923 23851
rect 19625 23817 19659 23851
rect 19993 23817 20027 23851
rect 22201 23817 22235 23851
rect 22661 23817 22695 23851
rect 23765 23817 23799 23851
rect 24777 23817 24811 23851
rect 30021 23817 30055 23851
rect 31217 23817 31251 23851
rect 32873 23817 32907 23851
rect 34805 23817 34839 23851
rect 22569 23749 22603 23783
rect 25973 23749 26007 23783
rect 28733 23749 28767 23783
rect 34437 23749 34471 23783
rect 17049 23681 17083 23715
rect 18705 23681 18739 23715
rect 20085 23681 20119 23715
rect 23489 23681 23523 23715
rect 23581 23681 23615 23715
rect 24593 23681 24627 23715
rect 28825 23681 28859 23715
rect 29837 23681 29871 23715
rect 30849 23681 30883 23715
rect 31033 23681 31067 23715
rect 32689 23681 32723 23715
rect 35265 23681 35299 23715
rect 35817 23681 35851 23715
rect 16773 23613 16807 23647
rect 16957 23613 16991 23647
rect 17969 23613 18003 23647
rect 20269 23613 20303 23647
rect 22845 23613 22879 23647
rect 26065 23613 26099 23647
rect 26157 23613 26191 23647
rect 27905 23613 27939 23647
rect 28917 23613 28951 23647
rect 29653 23613 29687 23647
rect 32505 23613 32539 23647
rect 33333 23613 33367 23647
rect 34161 23613 34195 23647
rect 34345 23613 34379 23647
rect 25605 23545 25639 23579
rect 26985 23545 27019 23579
rect 21189 23477 21223 23511
rect 28365 23477 28399 23511
rect 36461 23477 36495 23511
rect 17509 23273 17543 23307
rect 21097 23273 21131 23307
rect 24777 23273 24811 23307
rect 26617 23273 26651 23307
rect 29561 23273 29595 23307
rect 30205 23273 30239 23307
rect 31769 23273 31803 23307
rect 32505 23273 32539 23307
rect 34713 23273 34747 23307
rect 35541 23273 35575 23307
rect 36829 23273 36863 23307
rect 33333 23205 33367 23239
rect 19717 23137 19751 23171
rect 20545 23137 20579 23171
rect 22293 23137 22327 23171
rect 29009 23137 29043 23171
rect 33885 23137 33919 23171
rect 35081 23137 35115 23171
rect 35909 23137 35943 23171
rect 19901 23069 19935 23103
rect 20729 23069 20763 23103
rect 23029 23069 23063 23103
rect 23673 23069 23707 23103
rect 24501 23069 24535 23103
rect 24593 23069 24627 23103
rect 25237 23069 25271 23103
rect 28273 23069 28307 23103
rect 28457 23069 28491 23103
rect 30757 23069 30791 23103
rect 30941 23069 30975 23103
rect 31125 23069 31159 23103
rect 31585 23069 31619 23103
rect 32965 23069 32999 23103
rect 33149 23069 33183 23103
rect 34897 23069 34931 23103
rect 35725 23069 35759 23103
rect 37013 23069 37047 23103
rect 20637 23001 20671 23035
rect 21741 22933 21775 22967
rect 23121 22933 23155 22967
rect 25421 22933 25455 22967
rect 28089 22933 28123 22967
rect 23397 22729 23431 22763
rect 28549 22729 28583 22763
rect 30021 22729 30055 22763
rect 30757 22729 30791 22763
rect 32321 22729 32355 22763
rect 33333 22729 33367 22763
rect 33885 22729 33919 22763
rect 35265 22729 35299 22763
rect 35633 22729 35667 22763
rect 23857 22661 23891 22695
rect 24409 22661 24443 22695
rect 35725 22661 35759 22695
rect 20821 22593 20855 22627
rect 22201 22593 22235 22627
rect 23029 22593 23063 22627
rect 23213 22593 23247 22627
rect 25605 22593 25639 22627
rect 25789 22593 25823 22627
rect 27077 22593 27111 22627
rect 27721 22593 27755 22627
rect 28365 22593 28399 22627
rect 29837 22593 29871 22627
rect 32137 22593 32171 22627
rect 34069 22593 34103 22627
rect 21097 22525 21131 22559
rect 21925 22525 21959 22559
rect 22109 22525 22143 22559
rect 25421 22525 25455 22559
rect 29653 22525 29687 22559
rect 34253 22525 34287 22559
rect 35817 22525 35851 22559
rect 22569 22457 22603 22491
rect 27905 22457 27939 22491
rect 27261 22389 27295 22423
rect 34713 22389 34747 22423
rect 26157 22185 26191 22219
rect 28457 22185 28491 22219
rect 33425 22185 33459 22219
rect 34713 22185 34747 22219
rect 35909 22185 35943 22219
rect 23305 22117 23339 22151
rect 25605 22049 25639 22083
rect 26801 22049 26835 22083
rect 27629 22049 27663 22083
rect 28825 22049 28859 22083
rect 29837 22049 29871 22083
rect 30205 22049 30239 22083
rect 33977 22049 34011 22083
rect 35265 22049 35299 22083
rect 36461 22049 36495 22083
rect 21833 21981 21867 22015
rect 22753 21981 22787 22015
rect 27813 21981 27847 22015
rect 28641 21981 28675 22015
rect 30021 21981 30055 22015
rect 33793 21981 33827 22015
rect 35081 21981 35115 22015
rect 36277 21981 36311 22015
rect 26525 21913 26559 21947
rect 22109 21845 22143 21879
rect 26617 21845 26651 21879
rect 27997 21845 28031 21879
rect 33885 21845 33919 21879
rect 35173 21845 35207 21879
rect 36369 21845 36403 21879
rect 37197 21845 37231 21879
rect 28641 21641 28675 21675
rect 30849 21641 30883 21675
rect 31217 21641 31251 21675
rect 32781 21641 32815 21675
rect 36461 21641 36495 21675
rect 31309 21573 31343 21607
rect 32137 21573 32171 21607
rect 28273 21505 28307 21539
rect 30297 21505 30331 21539
rect 36277 21505 36311 21539
rect 28089 21437 28123 21471
rect 28181 21437 28215 21471
rect 31401 21437 31435 21471
rect 36093 21437 36127 21471
rect 27077 21301 27111 21335
rect 29193 21301 29227 21335
rect 29653 21301 29687 21335
rect 34253 21301 34287 21335
rect 35541 21301 35575 21335
rect 27261 21097 27295 21131
rect 27997 21097 28031 21131
rect 29745 21097 29779 21131
rect 30941 21097 30975 21131
rect 35725 21097 35759 21131
rect 36921 21097 36955 21131
rect 28549 20961 28583 20995
rect 30297 20961 30331 20995
rect 31493 20961 31527 20995
rect 36277 20961 36311 20995
rect 30113 20893 30147 20927
rect 31309 20893 31343 20927
rect 36093 20893 36127 20927
rect 28365 20825 28399 20859
rect 35265 20825 35299 20859
rect 36185 20825 36219 20859
rect 21005 20757 21039 20791
rect 28457 20757 28491 20791
rect 30205 20757 30239 20791
rect 31401 20757 31435 20791
rect 32229 20757 32263 20791
rect 20453 20553 20487 20587
rect 28365 20553 28399 20587
rect 29561 20553 29595 20587
rect 31309 20553 31343 20587
rect 20545 20417 20579 20451
rect 21833 20417 21867 20451
rect 29929 20417 29963 20451
rect 20729 20349 20763 20383
rect 30021 20349 30055 20383
rect 30205 20349 30239 20383
rect 20085 20213 20119 20247
rect 28825 20213 28859 20247
rect 30757 20213 30791 20247
rect 22845 20009 22879 20043
rect 29009 20009 29043 20043
rect 30481 20009 30515 20043
rect 36093 20009 36127 20043
rect 20453 19873 20487 19907
rect 21189 19873 21223 19907
rect 29561 19873 29595 19907
rect 35633 19873 35667 19907
rect 36645 19873 36679 19907
rect 21281 19805 21315 19839
rect 29745 19805 29779 19839
rect 36461 19805 36495 19839
rect 20177 19737 20211 19771
rect 22293 19737 22327 19771
rect 19809 19669 19843 19703
rect 20269 19669 20303 19703
rect 21373 19669 21407 19703
rect 21741 19669 21775 19703
rect 29929 19669 29963 19703
rect 36553 19669 36587 19703
rect 20453 19465 20487 19499
rect 21833 19465 21867 19499
rect 30297 19465 30331 19499
rect 35541 19465 35575 19499
rect 35909 19465 35943 19499
rect 20545 19329 20579 19363
rect 30113 19329 30147 19363
rect 21189 19261 21223 19295
rect 36001 19261 36035 19295
rect 29469 19125 29503 19159
rect 35081 19125 35115 19159
rect 35699 19125 35733 19159
rect 23581 18921 23615 18955
rect 36369 18921 36403 18955
rect 22385 18785 22419 18819
rect 22201 18717 22235 18751
rect 22109 18649 22143 18683
rect 23029 18649 23063 18683
rect 21741 18581 21775 18615
rect 17693 18377 17727 18411
rect 18521 18377 18555 18411
rect 33793 18377 33827 18411
rect 34253 18377 34287 18411
rect 17601 18241 17635 18275
rect 33885 18241 33919 18275
rect 34713 18241 34747 18275
rect 17877 18173 17911 18207
rect 33609 18173 33643 18207
rect 17233 18037 17267 18071
rect 33057 18037 33091 18071
rect 34897 18037 34931 18071
rect 34713 17833 34747 17867
rect 18061 17493 18095 17527
rect 19073 17289 19107 17323
rect 27077 17289 27111 17323
rect 25513 17153 25547 17187
rect 25237 17085 25271 17119
rect 25421 17085 25455 17119
rect 19533 17017 19567 17051
rect 25881 17017 25915 17051
rect 26341 16949 26375 16983
rect 22385 16745 22419 16779
rect 18429 16609 18463 16643
rect 18613 16609 18647 16643
rect 21005 16609 21039 16643
rect 21097 16609 21131 16643
rect 19717 16473 19751 16507
rect 17969 16405 18003 16439
rect 18337 16405 18371 16439
rect 20545 16405 20579 16439
rect 20913 16405 20947 16439
rect 21741 16405 21775 16439
rect 17417 16201 17451 16235
rect 19165 16201 19199 16235
rect 19073 16133 19107 16167
rect 19993 16133 20027 16167
rect 23213 16133 23247 16167
rect 24501 16133 24535 16167
rect 22017 16065 22051 16099
rect 23121 16065 23155 16099
rect 23949 16065 23983 16099
rect 18981 15997 19015 16031
rect 22201 15997 22235 16031
rect 23305 15997 23339 16031
rect 19533 15861 19567 15895
rect 21833 15861 21867 15895
rect 22753 15861 22787 15895
rect 21281 15657 21315 15691
rect 24593 15657 24627 15691
rect 21925 15589 21959 15623
rect 26617 15589 26651 15623
rect 16957 15521 16991 15555
rect 17141 15521 17175 15555
rect 20453 15521 20487 15555
rect 20637 15521 20671 15555
rect 36093 15521 36127 15555
rect 37105 15521 37139 15555
rect 17877 15453 17911 15487
rect 18061 15453 18095 15487
rect 21741 15453 21775 15487
rect 22385 15453 22419 15487
rect 22569 15453 22603 15487
rect 22753 15453 22787 15487
rect 23213 15453 23247 15487
rect 24409 15453 24443 15487
rect 26249 15453 26283 15487
rect 26453 15453 26487 15487
rect 27813 15453 27847 15487
rect 28365 15453 28399 15487
rect 37749 15453 37783 15487
rect 16865 15385 16899 15419
rect 16497 15317 16531 15351
rect 18245 15317 18279 15351
rect 19993 15317 20027 15351
rect 20361 15317 20395 15351
rect 23397 15317 23431 15351
rect 25421 15317 25455 15351
rect 36553 15317 36587 15351
rect 36921 15317 36955 15351
rect 37013 15317 37047 15351
rect 37933 15317 37967 15351
rect 18337 15113 18371 15147
rect 21833 15113 21867 15147
rect 23857 15113 23891 15147
rect 24961 15113 24995 15147
rect 32505 15113 32539 15147
rect 19901 15045 19935 15079
rect 22293 15045 22327 15079
rect 24869 15045 24903 15079
rect 19809 14977 19843 15011
rect 22201 14977 22235 15011
rect 23673 14977 23707 15011
rect 26249 14977 26283 15011
rect 30297 14977 30331 15011
rect 32137 14977 32171 15011
rect 32321 14977 32355 15011
rect 19993 14909 20027 14943
rect 22385 14909 22419 14943
rect 23489 14909 23523 14943
rect 25145 14909 25179 14943
rect 26065 14909 26099 14943
rect 20913 14841 20947 14875
rect 24501 14841 24535 14875
rect 31493 14841 31527 14875
rect 17233 14773 17267 14807
rect 17693 14773 17727 14807
rect 19441 14773 19475 14807
rect 26433 14773 26467 14807
rect 30481 14773 30515 14807
rect 19257 14569 19291 14603
rect 20545 14569 20579 14603
rect 21005 14569 21039 14603
rect 22661 14569 22695 14603
rect 25329 14569 25363 14603
rect 26433 14569 26467 14603
rect 25789 14501 25823 14535
rect 17233 14433 17267 14467
rect 18429 14433 18463 14467
rect 24777 14433 24811 14467
rect 36277 14433 36311 14467
rect 36461 14433 36495 14467
rect 15301 14365 15335 14399
rect 15485 14365 15519 14399
rect 28549 14365 28583 14399
rect 32413 14365 32447 14399
rect 32597 14365 32631 14399
rect 32781 14365 32815 14399
rect 33241 14365 33275 14399
rect 16957 14297 16991 14331
rect 24869 14297 24903 14331
rect 15669 14229 15703 14263
rect 16589 14229 16623 14263
rect 17049 14229 17083 14263
rect 17785 14229 17819 14263
rect 18153 14229 18187 14263
rect 18245 14229 18279 14263
rect 24961 14229 24995 14263
rect 28733 14229 28767 14263
rect 31861 14229 31895 14263
rect 33425 14229 33459 14263
rect 35633 14229 35667 14263
rect 36553 14229 36587 14263
rect 36921 14229 36955 14263
rect 16865 14025 16899 14059
rect 18705 14025 18739 14059
rect 25421 14025 25455 14059
rect 16681 13889 16715 13923
rect 17693 13889 17727 13923
rect 20177 13889 20211 13923
rect 20361 13889 20395 13923
rect 36461 13889 36495 13923
rect 15853 13821 15887 13855
rect 17509 13821 17543 13855
rect 17877 13821 17911 13855
rect 19993 13685 20027 13719
rect 36277 13685 36311 13719
rect 19441 13481 19475 13515
rect 36737 13481 36771 13515
rect 21649 13413 21683 13447
rect 24501 13413 24535 13447
rect 14381 13277 14415 13311
rect 15577 13277 15611 13311
rect 16129 13277 16163 13311
rect 16681 13277 16715 13311
rect 16773 13277 16807 13311
rect 18245 13277 18279 13311
rect 19257 13277 19291 13311
rect 19901 13277 19935 13311
rect 23029 13277 23063 13311
rect 25881 13277 25915 13311
rect 27721 13277 27755 13311
rect 32597 13277 32631 13311
rect 38117 13277 38151 13311
rect 22762 13209 22796 13243
rect 25614 13209 25648 13243
rect 27454 13209 27488 13243
rect 32330 13209 32364 13243
rect 37850 13209 37884 13243
rect 14565 13141 14599 13175
rect 16957 13141 16991 13175
rect 17509 13141 17543 13175
rect 18429 13141 18463 13175
rect 20085 13141 20119 13175
rect 26341 13141 26375 13175
rect 31217 13141 31251 13175
rect 32137 12937 32171 12971
rect 33977 12937 34011 12971
rect 37473 12937 37507 12971
rect 16129 12869 16163 12903
rect 30490 12869 30524 12903
rect 33272 12869 33306 12903
rect 15945 12801 15979 12835
rect 16865 12801 16899 12835
rect 17509 12801 17543 12835
rect 18981 12801 19015 12835
rect 19809 12801 19843 12835
rect 20637 12801 20671 12835
rect 22946 12801 22980 12835
rect 24786 12801 24820 12835
rect 25053 12801 25087 12835
rect 28650 12801 28684 12835
rect 28917 12801 28951 12835
rect 33517 12801 33551 12835
rect 35090 12801 35124 12835
rect 35357 12801 35391 12835
rect 37289 12801 37323 12835
rect 15301 12733 15335 12767
rect 15761 12733 15795 12767
rect 16681 12733 16715 12767
rect 18337 12733 18371 12767
rect 18797 12733 18831 12767
rect 19625 12733 19659 12767
rect 20821 12733 20855 12767
rect 23213 12733 23247 12767
rect 30757 12733 30791 12767
rect 17693 12665 17727 12699
rect 17049 12597 17083 12631
rect 19165 12597 19199 12631
rect 19993 12597 20027 12631
rect 20453 12597 20487 12631
rect 21833 12597 21867 12631
rect 23673 12597 23707 12631
rect 27537 12597 27571 12631
rect 29377 12597 29411 12631
rect 18337 12393 18371 12427
rect 20085 12393 20119 12427
rect 21649 12393 21683 12427
rect 25789 12393 25823 12427
rect 37473 12393 37507 12427
rect 15485 12257 15519 12291
rect 19625 12257 19659 12291
rect 27169 12257 27203 12291
rect 14933 12189 14967 12223
rect 15945 12189 15979 12223
rect 16129 12189 16163 12223
rect 17509 12189 17543 12223
rect 18153 12189 18187 12223
rect 19441 12189 19475 12223
rect 22762 12189 22796 12223
rect 23029 12189 23063 12223
rect 26902 12189 26936 12223
rect 29009 12189 29043 12223
rect 30858 12189 30892 12223
rect 31125 12189 31159 12223
rect 36093 12189 36127 12223
rect 16773 12121 16807 12155
rect 16957 12121 16991 12155
rect 28742 12121 28776 12155
rect 36360 12121 36394 12155
rect 16313 12053 16347 12087
rect 17693 12053 17727 12087
rect 19257 12053 19291 12087
rect 27629 12053 27663 12087
rect 29745 12053 29779 12087
rect 17509 11849 17543 11883
rect 18613 11849 18647 11883
rect 24133 11849 24167 11883
rect 32229 11849 32263 11883
rect 17049 11781 17083 11815
rect 20177 11781 20211 11815
rect 25246 11781 25280 11815
rect 33342 11781 33376 11815
rect 15577 11713 15611 11747
rect 17141 11713 17175 11747
rect 18521 11713 18555 11747
rect 19533 11713 19567 11747
rect 22946 11713 22980 11747
rect 25513 11713 25547 11747
rect 28190 11713 28224 11747
rect 28457 11713 28491 11747
rect 33609 11713 33643 11747
rect 16957 11645 16991 11679
rect 18705 11645 18739 11679
rect 23213 11645 23247 11679
rect 18153 11577 18187 11611
rect 15761 11509 15795 11543
rect 19717 11509 19751 11543
rect 21833 11509 21867 11543
rect 27077 11509 27111 11543
rect 14197 11305 14231 11339
rect 15485 11305 15519 11339
rect 17417 11305 17451 11339
rect 18061 11305 18095 11339
rect 30389 11305 30423 11339
rect 34713 11305 34747 11339
rect 36737 11305 36771 11339
rect 13553 11237 13587 11271
rect 16129 11237 16163 11271
rect 16773 11237 16807 11271
rect 18705 11237 18739 11271
rect 14657 11169 14691 11203
rect 14841 11169 14875 11203
rect 26617 11169 26651 11203
rect 38117 11169 38151 11203
rect 13369 11101 13403 11135
rect 15945 11101 15979 11135
rect 16589 11101 16623 11135
rect 17233 11101 17267 11135
rect 17877 11101 17911 11135
rect 18521 11101 18555 11135
rect 19257 11101 19291 11135
rect 23121 11101 23155 11135
rect 31502 11101 31536 11135
rect 31769 11101 31803 11135
rect 32229 11101 32263 11135
rect 36093 11101 36127 11135
rect 14565 11033 14599 11067
rect 22854 11033 22888 11067
rect 26350 11033 26384 11067
rect 32474 11033 32508 11067
rect 35826 11033 35860 11067
rect 37850 11033 37884 11067
rect 19441 10965 19475 10999
rect 21741 10965 21775 10999
rect 25237 10965 25271 10999
rect 33609 10965 33643 10999
rect 15853 10761 15887 10795
rect 19441 10761 19475 10795
rect 15393 10693 15427 10727
rect 16773 10693 16807 10727
rect 35541 10693 35575 10727
rect 11529 10625 11563 10659
rect 15485 10625 15519 10659
rect 18061 10625 18095 10659
rect 19349 10625 19383 10659
rect 20085 10625 20119 10659
rect 25145 10625 25179 10659
rect 28549 10625 28583 10659
rect 28805 10625 28839 10659
rect 33793 10625 33827 10659
rect 15301 10557 15335 10591
rect 18797 10557 18831 10591
rect 11713 10489 11747 10523
rect 18245 10489 18279 10523
rect 23857 10489 23891 10523
rect 20269 10421 20303 10455
rect 29929 10421 29963 10455
rect 38025 10421 38059 10455
rect 15945 10217 15979 10251
rect 16497 10217 16531 10251
rect 18337 10217 18371 10251
rect 27353 10217 27387 10251
rect 15393 10081 15427 10115
rect 15485 10081 15519 10115
rect 17785 10081 17819 10115
rect 23213 10081 23247 10115
rect 19809 10013 19843 10047
rect 19901 10013 19935 10047
rect 20085 10013 20119 10047
rect 20545 10013 20579 10047
rect 26065 10013 26099 10047
rect 31217 10013 31251 10047
rect 15577 9945 15611 9979
rect 17877 9945 17911 9979
rect 22946 9945 22980 9979
rect 17969 9877 18003 9911
rect 20729 9877 20763 9911
rect 21833 9877 21867 9911
rect 32505 9877 32539 9911
rect 37381 9877 37415 9911
rect 37841 9877 37875 9911
rect 11529 9673 11563 9707
rect 18521 9673 18555 9707
rect 20913 9673 20947 9707
rect 10793 9605 10827 9639
rect 11989 9605 12023 9639
rect 14381 9605 14415 9639
rect 15209 9605 15243 9639
rect 25154 9605 25188 9639
rect 30398 9605 30432 9639
rect 34170 9605 34204 9639
rect 11897 9537 11931 9571
rect 14289 9537 14323 9571
rect 16865 9537 16899 9571
rect 19073 9537 19107 9571
rect 19257 9537 19291 9571
rect 19441 9537 19475 9571
rect 20085 9537 20119 9571
rect 20729 9537 20763 9571
rect 22201 9537 22235 9571
rect 22457 9537 22491 9571
rect 25421 9537 25455 9571
rect 28098 9537 28132 9571
rect 28365 9537 28399 9571
rect 30665 9537 30699 9571
rect 34437 9537 34471 9571
rect 34897 9537 34931 9571
rect 35153 9537 35187 9571
rect 12081 9469 12115 9503
rect 12817 9469 12851 9503
rect 14565 9469 14599 9503
rect 16773 9469 16807 9503
rect 13921 9401 13955 9435
rect 20269 9401 20303 9435
rect 23581 9401 23615 9435
rect 16037 9333 16071 9367
rect 17233 9333 17267 9367
rect 17785 9333 17819 9367
rect 24041 9333 24075 9367
rect 26985 9333 27019 9367
rect 29285 9333 29319 9367
rect 33057 9333 33091 9367
rect 36277 9333 36311 9367
rect 37749 9333 37783 9367
rect 14289 9129 14323 9163
rect 18705 9129 18739 9163
rect 19993 9129 20027 9163
rect 26433 9129 26467 9163
rect 27445 9129 27479 9163
rect 30573 9129 30607 9163
rect 33241 9129 33275 9163
rect 34897 9129 34931 9163
rect 14841 9061 14875 9095
rect 17509 9061 17543 9095
rect 35633 9061 35667 9095
rect 10057 8993 10091 9027
rect 10241 8993 10275 9027
rect 16957 8993 16991 9027
rect 19349 8993 19383 9027
rect 19533 8993 19567 9027
rect 20545 8993 20579 9027
rect 22937 8993 22971 9027
rect 11621 8925 11655 8959
rect 12265 8925 12299 8959
rect 14105 8925 14139 8959
rect 17509 8925 17543 8959
rect 17693 8925 17727 8959
rect 25078 8925 25112 8959
rect 28825 8925 28859 8959
rect 31686 8925 31720 8959
rect 31953 8925 31987 8959
rect 34713 8925 34747 8959
rect 37013 8925 37047 8959
rect 10333 8857 10367 8891
rect 22670 8857 22704 8891
rect 25298 8857 25332 8891
rect 28558 8857 28592 8891
rect 36746 8857 36780 8891
rect 10701 8789 10735 8823
rect 11713 8789 11747 8823
rect 19625 8789 19659 8823
rect 21005 8789 21039 8823
rect 21557 8789 21591 8823
rect 33885 8789 33919 8823
rect 37473 8789 37507 8823
rect 38025 8789 38059 8823
rect 10885 8585 10919 8619
rect 11989 8585 12023 8619
rect 13921 8585 13955 8619
rect 14381 8585 14415 8619
rect 15945 8585 15979 8619
rect 34161 8585 34195 8619
rect 36277 8585 36311 8619
rect 12081 8517 12115 8551
rect 20453 8517 20487 8551
rect 21005 8517 21039 8551
rect 35817 8517 35851 8551
rect 10701 8449 10735 8483
rect 13185 8449 13219 8483
rect 14289 8449 14323 8483
rect 15209 8449 15243 8483
rect 15393 8449 15427 8483
rect 18061 8449 18095 8483
rect 18613 8449 18647 8483
rect 22946 8449 22980 8483
rect 23213 8449 23247 8483
rect 28098 8449 28132 8483
rect 28365 8449 28399 8483
rect 33977 8449 34011 8483
rect 11897 8381 11931 8415
rect 14565 8381 14599 8415
rect 19809 8381 19843 8415
rect 20177 8381 20211 8415
rect 20269 8381 20303 8415
rect 12449 8313 12483 8347
rect 13369 8313 13403 8347
rect 21833 8313 21867 8347
rect 26985 8313 27019 8347
rect 37381 8313 37415 8347
rect 37933 8313 37967 8347
rect 15301 8245 15335 8279
rect 32229 8245 32263 8279
rect 33333 8245 33367 8279
rect 34621 8245 34655 8279
rect 35173 8245 35207 8279
rect 11069 8041 11103 8075
rect 12633 8041 12667 8075
rect 18061 8041 18095 8075
rect 30481 8041 30515 8075
rect 34713 8041 34747 8075
rect 38117 8041 38151 8075
rect 18705 7973 18739 8007
rect 16589 7905 16623 7939
rect 19901 7905 19935 7939
rect 32413 7905 32447 7939
rect 35173 7905 35207 7939
rect 35357 7905 35391 7939
rect 15209 7837 15243 7871
rect 15393 7837 15427 7871
rect 15945 7837 15979 7871
rect 17877 7837 17911 7871
rect 18521 7837 18555 7871
rect 19257 7837 19291 7871
rect 23121 7837 23155 7871
rect 27629 7837 27663 7871
rect 31953 7837 31987 7871
rect 36093 7837 36127 7871
rect 36737 7837 36771 7871
rect 22854 7769 22888 7803
rect 27362 7769 27396 7803
rect 32658 7769 32692 7803
rect 36993 7769 37027 7803
rect 16037 7701 16071 7735
rect 19441 7701 19475 7735
rect 21741 7701 21775 7735
rect 26249 7701 26283 7735
rect 33793 7701 33827 7735
rect 35081 7701 35115 7735
rect 36277 7701 36311 7735
rect 10517 7497 10551 7531
rect 12081 7497 12115 7531
rect 15577 7497 15611 7531
rect 16037 7497 16071 7531
rect 16957 7497 16991 7531
rect 17417 7497 17451 7531
rect 18705 7497 18739 7531
rect 19625 7497 19659 7531
rect 20177 7497 20211 7531
rect 29101 7497 29135 7531
rect 29561 7497 29595 7531
rect 34805 7497 34839 7531
rect 35357 7497 35391 7531
rect 10609 7429 10643 7463
rect 24286 7429 24320 7463
rect 30674 7429 30708 7463
rect 34345 7429 34379 7463
rect 36461 7429 36495 7463
rect 9597 7361 9631 7395
rect 11897 7361 11931 7395
rect 13553 7361 13587 7395
rect 13737 7361 13771 7395
rect 15209 7361 15243 7395
rect 15393 7361 15427 7395
rect 17049 7361 17083 7395
rect 18337 7361 18371 7395
rect 19441 7361 19475 7395
rect 28917 7361 28951 7395
rect 32137 7361 32171 7395
rect 34437 7361 34471 7395
rect 10425 7293 10459 7327
rect 14197 7293 14231 7327
rect 16773 7293 16807 7327
rect 18153 7293 18187 7327
rect 18245 7293 18279 7327
rect 24041 7293 24075 7327
rect 30941 7293 30975 7327
rect 34161 7293 34195 7327
rect 37841 7293 37875 7327
rect 9781 7225 9815 7259
rect 35817 7225 35851 7259
rect 37289 7225 37323 7259
rect 10977 7157 11011 7191
rect 13001 7157 13035 7191
rect 13645 7157 13679 7191
rect 25421 7157 25455 7191
rect 31401 7157 31435 7191
rect 32321 7157 32355 7191
rect 32781 7157 32815 7191
rect 33609 7157 33643 7191
rect 15945 6953 15979 6987
rect 17877 6953 17911 6987
rect 19257 6953 19291 6987
rect 31677 6885 31711 6919
rect 12541 6817 12575 6851
rect 14289 6817 14323 6851
rect 14473 6817 14507 6851
rect 15393 6817 15427 6851
rect 16405 6817 16439 6851
rect 18705 6817 18739 6851
rect 19809 6817 19843 6851
rect 30573 6817 30607 6851
rect 30757 6817 30791 6851
rect 35173 6817 35207 6851
rect 35357 6817 35391 6851
rect 36185 6817 36219 6851
rect 11529 6749 11563 6783
rect 13093 6749 13127 6783
rect 14381 6749 14415 6783
rect 14565 6749 14599 6783
rect 16589 6749 16623 6783
rect 16773 6749 16807 6783
rect 17233 6749 17267 6783
rect 20453 6749 20487 6783
rect 23029 6749 23063 6783
rect 26902 6749 26936 6783
rect 27169 6749 27203 6783
rect 33057 6749 33091 6783
rect 33977 6749 34011 6783
rect 35081 6749 35115 6783
rect 13369 6681 13403 6715
rect 22762 6681 22796 6715
rect 29929 6681 29963 6715
rect 32790 6681 32824 6715
rect 36430 6681 36464 6715
rect 38025 6681 38059 6715
rect 11069 6613 11103 6647
rect 11713 6613 11747 6647
rect 14105 6613 14139 6647
rect 17417 6613 17451 6647
rect 19625 6613 19659 6647
rect 19717 6613 19751 6647
rect 20637 6613 20671 6647
rect 21649 6613 21683 6647
rect 25789 6613 25823 6647
rect 30849 6613 30883 6647
rect 31217 6613 31251 6647
rect 34161 6613 34195 6647
rect 34713 6613 34747 6647
rect 37565 6613 37599 6647
rect 9965 6409 9999 6443
rect 11897 6409 11931 6443
rect 12265 6409 12299 6443
rect 13921 6409 13955 6443
rect 18981 6409 19015 6443
rect 19441 6409 19475 6443
rect 20177 6409 20211 6443
rect 28457 6409 28491 6443
rect 30297 6409 30331 6443
rect 30757 6409 30791 6443
rect 32413 6409 32447 6443
rect 32873 6409 32907 6443
rect 35817 6409 35851 6443
rect 10517 6341 10551 6375
rect 11805 6341 11839 6375
rect 14749 6341 14783 6375
rect 15117 6341 15151 6375
rect 18337 6341 18371 6375
rect 24746 6341 24780 6375
rect 31493 6341 31527 6375
rect 10885 6273 10919 6307
rect 12725 6273 12759 6307
rect 12909 6273 12943 6307
rect 13553 6273 13587 6307
rect 13737 6273 13771 6307
rect 15761 6273 15795 6307
rect 16129 6273 16163 6307
rect 16773 6273 16807 6307
rect 18245 6273 18279 6307
rect 18429 6273 18463 6307
rect 22946 6273 22980 6307
rect 29570 6273 29604 6307
rect 29837 6273 29871 6307
rect 30665 6273 30699 6307
rect 32505 6273 32539 6307
rect 34621 6273 34655 6307
rect 37657 6273 37691 6307
rect 11621 6205 11655 6239
rect 16957 6205 16991 6239
rect 23213 6205 23247 6239
rect 24501 6205 24535 6239
rect 30849 6205 30883 6239
rect 32321 6205 32355 6239
rect 21097 6137 21131 6171
rect 33885 6137 33919 6171
rect 12725 6069 12759 6103
rect 15577 6069 15611 6103
rect 15761 6069 15795 6103
rect 17693 6069 17727 6103
rect 21833 6069 21867 6103
rect 25881 6069 25915 6103
rect 33333 6069 33367 6103
rect 34805 6069 34839 6103
rect 35357 6069 35391 6103
rect 36369 6069 36403 6103
rect 37473 6069 37507 6103
rect 9965 5865 9999 5899
rect 12081 5865 12115 5899
rect 12909 5865 12943 5899
rect 15485 5865 15519 5899
rect 17325 5865 17359 5899
rect 26893 5865 26927 5899
rect 29561 5865 29595 5899
rect 31401 5865 31435 5899
rect 33609 5865 33643 5899
rect 34713 5865 34747 5899
rect 36001 5865 36035 5899
rect 38117 5865 38151 5899
rect 11069 5797 11103 5831
rect 20545 5797 20579 5831
rect 22109 5797 22143 5831
rect 29009 5797 29043 5831
rect 32045 5797 32079 5831
rect 9413 5729 9447 5763
rect 9505 5729 9539 5763
rect 13369 5729 13403 5763
rect 16037 5729 16071 5763
rect 16681 5729 16715 5763
rect 18705 5729 18739 5763
rect 21373 5729 21407 5763
rect 35173 5729 35207 5763
rect 35357 5729 35391 5763
rect 36737 5729 36771 5763
rect 10885 5661 10919 5695
rect 12633 5661 12667 5695
rect 12909 5661 12943 5695
rect 14933 5661 14967 5695
rect 18153 5661 18187 5695
rect 20821 5661 20855 5695
rect 21281 5661 21315 5695
rect 21465 5661 21499 5695
rect 23222 5661 23256 5695
rect 23489 5661 23523 5695
rect 28006 5661 28040 5695
rect 28273 5661 28307 5695
rect 30941 5661 30975 5695
rect 36185 5661 36219 5695
rect 9597 5593 9631 5627
rect 11621 5593 11655 5627
rect 16957 5593 16991 5627
rect 17969 5593 18003 5627
rect 19717 5593 19751 5627
rect 20545 5593 20579 5627
rect 24869 5593 24903 5627
rect 30674 5593 30708 5627
rect 33057 5593 33091 5627
rect 36982 5593 37016 5627
rect 7941 5525 7975 5559
rect 12725 5525 12759 5559
rect 14381 5525 14415 5559
rect 16865 5525 16899 5559
rect 17785 5525 17819 5559
rect 19809 5525 19843 5559
rect 20729 5525 20763 5559
rect 32505 5525 32539 5559
rect 35081 5525 35115 5559
rect 8677 5321 8711 5355
rect 10517 5321 10551 5355
rect 10977 5321 11011 5355
rect 15669 5321 15703 5355
rect 19073 5321 19107 5355
rect 20361 5321 20395 5355
rect 36645 5321 36679 5355
rect 37933 5321 37967 5355
rect 15117 5253 15151 5287
rect 20177 5253 20211 5287
rect 25605 5253 25639 5287
rect 26249 5253 26283 5287
rect 28098 5253 28132 5287
rect 32873 5253 32907 5287
rect 33793 5253 33827 5287
rect 35541 5253 35575 5287
rect 10609 5185 10643 5219
rect 11529 5185 11563 5219
rect 11713 5185 11747 5219
rect 12909 5185 12943 5219
rect 13737 5185 13771 5219
rect 14013 5185 14047 5219
rect 14197 5185 14231 5219
rect 14841 5185 14875 5219
rect 15577 5185 15611 5219
rect 15853 5185 15887 5219
rect 16865 5185 16899 5219
rect 18061 5185 18095 5219
rect 18889 5185 18923 5219
rect 19993 5185 20027 5219
rect 21005 5185 21039 5219
rect 25145 5185 25179 5219
rect 36001 5185 36035 5219
rect 37473 5185 37507 5219
rect 38117 5185 38151 5219
rect 10425 5117 10459 5151
rect 12633 5117 12667 5151
rect 13875 5117 13909 5151
rect 14933 5117 14967 5151
rect 17049 5117 17083 5151
rect 17141 5117 17175 5151
rect 23489 5117 23523 5151
rect 28365 5117 28399 5151
rect 32597 5117 32631 5151
rect 32781 5117 32815 5151
rect 9229 5049 9263 5083
rect 12725 5049 12759 5083
rect 16681 5049 16715 5083
rect 20913 5049 20947 5083
rect 26985 5049 27019 5083
rect 33241 5049 33275 5083
rect 37289 5049 37323 5083
rect 7573 4981 7607 5015
rect 8125 4981 8159 5015
rect 9781 4981 9815 5015
rect 11897 4981 11931 5015
rect 13093 4981 13127 5015
rect 14105 4981 14139 5015
rect 14657 4981 14691 5015
rect 15117 4981 15151 5015
rect 15853 4981 15887 5015
rect 18245 4981 18279 5015
rect 21833 4981 21867 5015
rect 28825 4981 28859 5015
rect 29377 4981 29411 5015
rect 29929 4981 29963 5015
rect 30573 4981 30607 5015
rect 31585 4981 31619 5015
rect 36185 4981 36219 5015
rect 11713 4777 11747 4811
rect 14473 4777 14507 4811
rect 16497 4777 16531 4811
rect 17141 4777 17175 4811
rect 17693 4777 17727 4811
rect 20361 4777 20395 4811
rect 21005 4777 21039 4811
rect 27077 4777 27111 4811
rect 31861 4777 31895 4811
rect 34161 4777 34195 4811
rect 35449 4777 35483 4811
rect 9413 4709 9447 4743
rect 10609 4709 10643 4743
rect 25237 4709 25271 4743
rect 37381 4709 37415 4743
rect 7849 4641 7883 4675
rect 30665 4641 30699 4675
rect 31217 4641 31251 4675
rect 34805 4641 34839 4675
rect 34989 4641 35023 4675
rect 7297 4573 7331 4607
rect 10425 4573 10459 4607
rect 12725 4573 12759 4607
rect 12909 4573 12943 4607
rect 13093 4573 13127 4607
rect 14197 4573 14231 4607
rect 14381 4573 14415 4607
rect 14473 4573 14507 4607
rect 15393 4573 15427 4607
rect 16589 4573 16623 4607
rect 18153 4573 18187 4607
rect 19533 4573 19567 4607
rect 23029 4573 23063 4607
rect 24593 4573 24627 4607
rect 26350 4573 26384 4607
rect 26617 4573 26651 4607
rect 28457 4573 28491 4607
rect 30113 4573 30147 4607
rect 32505 4573 32539 4607
rect 32965 4573 32999 4607
rect 33977 4573 34011 4607
rect 36001 4573 36035 4607
rect 36268 4573 36302 4607
rect 38117 4573 38151 4607
rect 6745 4505 6779 4539
rect 8401 4505 8435 4539
rect 11161 4505 11195 4539
rect 22762 4505 22796 4539
rect 23673 4505 23707 4539
rect 28190 4505 28224 4539
rect 31401 4505 31435 4539
rect 31493 4505 31527 4539
rect 5273 4437 5307 4471
rect 5917 4437 5951 4471
rect 9965 4437 9999 4471
rect 12265 4437 12299 4471
rect 15853 4437 15887 4471
rect 18337 4437 18371 4471
rect 19717 4437 19751 4471
rect 21649 4437 21683 4471
rect 24777 4437 24811 4471
rect 29009 4437 29043 4471
rect 29929 4437 29963 4471
rect 32321 4437 32355 4471
rect 33149 4437 33183 4471
rect 35081 4437 35115 4471
rect 37933 4437 37967 4471
rect 8309 4233 8343 4267
rect 10609 4233 10643 4267
rect 28457 4233 28491 4267
rect 28917 4233 28951 4267
rect 31493 4233 31527 4267
rect 32137 4233 32171 4267
rect 33793 4233 33827 4267
rect 34805 4233 34839 4267
rect 35357 4233 35391 4267
rect 19717 4165 19751 4199
rect 29828 4165 29862 4199
rect 32505 4165 32539 4199
rect 7757 4097 7791 4131
rect 10241 4097 10275 4131
rect 12081 4097 12115 4131
rect 12725 4097 12759 4131
rect 13369 4097 13403 4131
rect 13553 4097 13587 4131
rect 14013 4097 14047 4131
rect 15669 4097 15703 4131
rect 17233 4097 17267 4131
rect 17601 4097 17635 4131
rect 17785 4097 17819 4131
rect 18061 4097 18095 4131
rect 18245 4097 18279 4131
rect 18705 4097 18739 4131
rect 19625 4097 19659 4131
rect 20545 4097 20579 4131
rect 21189 4097 21223 4131
rect 22937 4097 22971 4131
rect 24133 4097 24167 4131
rect 24389 4097 24423 4131
rect 27333 4097 27367 4131
rect 29101 4097 29135 4131
rect 32597 4097 32631 4131
rect 34621 4097 34655 4131
rect 36470 4097 36504 4131
rect 36737 4097 36771 4131
rect 37473 4097 37507 4131
rect 38117 4097 38151 4131
rect 6653 4029 6687 4063
rect 10057 4029 10091 4063
rect 10149 4029 10183 4063
rect 11621 4029 11655 4063
rect 19441 4029 19475 4063
rect 27077 4029 27111 4063
rect 29561 4029 29595 4063
rect 32689 4029 32723 4063
rect 33517 4029 33551 4063
rect 33701 4029 33735 4063
rect 5825 3961 5859 3995
rect 8861 3961 8895 3995
rect 13369 3961 13403 3995
rect 15209 3961 15243 3995
rect 20085 3961 20119 3995
rect 21833 3961 21867 3995
rect 26065 3961 26099 3995
rect 30941 3961 30975 3995
rect 34161 3961 34195 3995
rect 37933 3961 37967 3995
rect 3985 3893 4019 3927
rect 4629 3893 4663 3927
rect 5273 3893 5307 3927
rect 7205 3893 7239 3927
rect 9413 3893 9447 3927
rect 12265 3893 12299 3927
rect 12909 3893 12943 3927
rect 14197 3893 14231 3927
rect 15853 3893 15887 3927
rect 16773 3893 16807 3927
rect 20729 3893 20763 3927
rect 22477 3893 22511 3927
rect 23489 3893 23523 3927
rect 25513 3893 25547 3927
rect 37289 3893 37323 3927
rect 7849 3689 7883 3723
rect 8401 3689 8435 3723
rect 10333 3689 10367 3723
rect 11713 3689 11747 3723
rect 14381 3689 14415 3723
rect 16681 3689 16715 3723
rect 18337 3689 18371 3723
rect 19257 3689 19291 3723
rect 22753 3689 22787 3723
rect 26525 3689 26559 3723
rect 29009 3689 29043 3723
rect 30113 3689 30147 3723
rect 36829 3689 36863 3723
rect 6193 3621 6227 3655
rect 7297 3621 7331 3655
rect 14657 3621 14691 3655
rect 15301 3621 15335 3655
rect 15393 3621 15427 3655
rect 28273 3621 28307 3655
rect 34989 3621 35023 3655
rect 6745 3553 6779 3587
rect 12173 3553 12207 3587
rect 14381 3553 14415 3587
rect 16497 3553 16531 3587
rect 17693 3553 17727 3587
rect 19717 3553 19751 3587
rect 19901 3553 19935 3587
rect 33517 3553 33551 3587
rect 36369 3553 36403 3587
rect 4077 3485 4111 3519
rect 5641 3485 5675 3519
rect 9137 3485 9171 3519
rect 10149 3485 10183 3519
rect 10885 3485 10919 3519
rect 11529 3485 11563 3519
rect 12424 3485 12458 3519
rect 12541 3485 12575 3519
rect 12633 3485 12667 3519
rect 13369 3485 13403 3519
rect 13553 3485 13587 3519
rect 14473 3485 14507 3519
rect 15393 3485 15427 3519
rect 16405 3485 16439 3519
rect 17877 3485 17911 3519
rect 20729 3485 20763 3519
rect 21373 3485 21407 3519
rect 21629 3485 21663 3519
rect 23489 3485 23523 3519
rect 24685 3485 24719 3519
rect 25421 3485 25455 3519
rect 27813 3485 27847 3519
rect 28457 3485 28491 3519
rect 29561 3485 29595 3519
rect 32965 3485 32999 3519
rect 37013 3485 37047 3519
rect 37657 3485 37691 3519
rect 5089 3417 5123 3451
rect 12311 3417 12345 3451
rect 13461 3417 13495 3451
rect 14197 3417 14231 3451
rect 15117 3417 15151 3451
rect 16681 3417 16715 3451
rect 17969 3417 18003 3451
rect 36124 3417 36158 3451
rect 3157 3349 3191 3383
rect 4261 3349 4295 3383
rect 9321 3349 9355 3383
rect 11069 3349 11103 3383
rect 12817 3349 12851 3383
rect 16221 3349 16255 3383
rect 19625 3349 19659 3383
rect 20545 3349 20579 3383
rect 23305 3349 23339 3383
rect 24501 3349 24535 3383
rect 25237 3349 25271 3383
rect 30665 3349 30699 3383
rect 31493 3349 31527 3383
rect 33701 3349 33735 3383
rect 33793 3349 33827 3383
rect 34161 3349 34195 3383
rect 37473 3349 37507 3383
rect 5825 3145 5859 3179
rect 7021 3145 7055 3179
rect 7757 3145 7791 3179
rect 9229 3145 9263 3179
rect 9597 3145 9631 3179
rect 14013 3145 14047 3179
rect 15577 3145 15611 3179
rect 15945 3145 15979 3179
rect 17417 3145 17451 3179
rect 17877 3145 17911 3179
rect 19993 3145 20027 3179
rect 23213 3145 23247 3179
rect 25881 3145 25915 3179
rect 28825 3145 28859 3179
rect 30849 3145 30883 3179
rect 31585 3145 31619 3179
rect 33977 3145 34011 3179
rect 35081 3145 35115 3179
rect 3065 3077 3099 3111
rect 26433 3077 26467 3111
rect 28098 3077 28132 3111
rect 29960 3077 29994 3111
rect 36216 3077 36250 3111
rect 38025 3077 38059 3111
rect 3801 3009 3835 3043
rect 4353 3009 4387 3043
rect 4997 3009 5031 3043
rect 5641 3009 5675 3043
rect 6837 3009 6871 3043
rect 7573 3009 7607 3043
rect 8217 3009 8251 3043
rect 10241 3009 10275 3043
rect 11989 3009 12023 3043
rect 13001 3009 13035 3043
rect 13645 3009 13679 3043
rect 14565 3009 14599 3043
rect 16957 3009 16991 3043
rect 17049 3009 17083 3043
rect 18153 3009 18187 3043
rect 18429 3009 18463 3043
rect 19625 3009 19659 3043
rect 20913 3009 20947 3043
rect 21833 3009 21867 3043
rect 22100 3009 22134 3043
rect 23949 3009 23983 3043
rect 24501 3009 24535 3043
rect 24757 3009 24791 3043
rect 28365 3009 28399 3043
rect 30665 3009 30699 3043
rect 31401 3009 31435 3043
rect 32393 3009 32427 3043
rect 34161 3009 34195 3043
rect 36461 3009 36495 3043
rect 9045 2941 9079 2975
rect 9137 2941 9171 2975
rect 10333 2941 10367 2975
rect 10609 2941 10643 2975
rect 11713 2941 11747 2975
rect 11897 2941 11931 2975
rect 13737 2941 13771 2975
rect 15301 2941 15335 2975
rect 15485 2941 15519 2975
rect 16865 2941 16899 2975
rect 19441 2941 19475 2975
rect 19533 2941 19567 2975
rect 30205 2941 30239 2975
rect 32137 2941 32171 2975
rect 4537 2873 4571 2907
rect 13185 2873 13219 2907
rect 23765 2873 23799 2907
rect 26985 2873 27019 2907
rect 1777 2805 1811 2839
rect 2329 2805 2363 2839
rect 3617 2805 3651 2839
rect 5181 2805 5215 2839
rect 8401 2805 8435 2839
rect 12357 2805 12391 2839
rect 13645 2805 13679 2839
rect 14749 2805 14783 2839
rect 18337 2805 18371 2839
rect 20729 2805 20763 2839
rect 33517 2805 33551 2839
rect 37933 2805 37967 2839
rect 7757 2601 7791 2635
rect 9873 2601 9907 2635
rect 10701 2601 10735 2635
rect 14841 2601 14875 2635
rect 16129 2601 16163 2635
rect 17141 2601 17175 2635
rect 19993 2601 20027 2635
rect 20453 2601 20487 2635
rect 28549 2601 28583 2635
rect 30849 2601 30883 2635
rect 33977 2601 34011 2635
rect 7113 2533 7147 2567
rect 8401 2533 8435 2567
rect 9229 2533 9263 2567
rect 22293 2533 22327 2567
rect 25973 2533 26007 2567
rect 27077 2533 27111 2567
rect 30389 2533 30423 2567
rect 35357 2533 35391 2567
rect 4077 2465 4111 2499
rect 10333 2465 10367 2499
rect 19349 2465 19383 2499
rect 23673 2465 23707 2499
rect 32597 2465 32631 2499
rect 36737 2465 36771 2499
rect 37565 2465 37599 2499
rect 1685 2397 1719 2431
rect 2421 2397 2455 2431
rect 2697 2397 2731 2431
rect 3801 2397 3835 2431
rect 5641 2397 5675 2431
rect 6929 2397 6963 2431
rect 7573 2397 7607 2431
rect 8217 2397 8251 2431
rect 9045 2397 9079 2431
rect 9689 2397 9723 2431
rect 10517 2397 10551 2431
rect 12081 2397 12115 2431
rect 12725 2397 12759 2431
rect 13369 2397 13403 2431
rect 14657 2397 14691 2431
rect 15301 2397 15335 2431
rect 16957 2397 16991 2431
rect 17693 2397 17727 2431
rect 18429 2397 18463 2431
rect 19533 2397 19567 2431
rect 21281 2397 21315 2431
rect 24685 2397 24719 2431
rect 25421 2397 25455 2431
rect 26157 2397 26191 2431
rect 27261 2397 27295 2431
rect 27997 2397 28031 2431
rect 28733 2397 28767 2431
rect 29745 2397 29779 2431
rect 30205 2397 30239 2431
rect 31033 2397 31067 2431
rect 31585 2397 31619 2431
rect 34897 2397 34931 2431
rect 36481 2397 36515 2431
rect 37289 2397 37323 2431
rect 19625 2329 19659 2363
rect 23406 2329 23440 2363
rect 32864 2329 32898 2363
rect 1869 2261 1903 2295
rect 5181 2261 5215 2295
rect 5825 2261 5859 2295
rect 6469 2261 6503 2295
rect 11621 2261 11655 2295
rect 12265 2261 12299 2295
rect 12909 2261 12943 2295
rect 13553 2261 13587 2295
rect 14197 2261 14231 2295
rect 15485 2261 15519 2295
rect 17877 2261 17911 2295
rect 18613 2261 18647 2295
rect 21097 2261 21131 2295
rect 24501 2261 24535 2295
rect 25237 2261 25271 2295
rect 27813 2261 27847 2295
rect 29561 2261 29595 2295
rect 34713 2261 34747 2295
<< metal1 >>
rect 21266 37680 21272 37732
rect 21324 37720 21330 37732
rect 23842 37720 23848 37732
rect 21324 37692 23848 37720
rect 21324 37680 21330 37692
rect 23842 37680 23848 37692
rect 23900 37680 23906 37732
rect 13446 37612 13452 37664
rect 13504 37652 13510 37664
rect 26234 37652 26240 37664
rect 13504 37624 26240 37652
rect 13504 37612 13510 37624
rect 26234 37612 26240 37624
rect 26292 37612 26298 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 20441 37451 20499 37457
rect 20441 37417 20453 37451
rect 20487 37448 20499 37451
rect 23842 37448 23848 37460
rect 20487 37420 22094 37448
rect 23755 37420 23848 37448
rect 20487 37417 20499 37420
rect 20441 37411 20499 37417
rect 1765 37383 1823 37389
rect 1765 37349 1777 37383
rect 1811 37380 1823 37383
rect 9950 37380 9956 37392
rect 1811 37352 9956 37380
rect 1811 37349 1823 37352
rect 1765 37343 1823 37349
rect 9950 37340 9956 37352
rect 10008 37340 10014 37392
rect 22066 37380 22094 37420
rect 23842 37408 23848 37420
rect 23900 37448 23906 37460
rect 28442 37448 28448 37460
rect 23900 37420 28448 37448
rect 23900 37408 23906 37420
rect 28442 37408 28448 37420
rect 28500 37408 28506 37460
rect 29362 37408 29368 37460
rect 29420 37448 29426 37460
rect 30377 37451 30435 37457
rect 30377 37448 30389 37451
rect 29420 37420 30389 37448
rect 29420 37408 29426 37420
rect 30377 37417 30389 37420
rect 30423 37417 30435 37451
rect 30377 37411 30435 37417
rect 35066 37380 35072 37392
rect 22066 37352 35072 37380
rect 35066 37340 35072 37352
rect 35124 37340 35130 37392
rect 17770 37272 17776 37324
rect 17828 37312 17834 37324
rect 17865 37315 17923 37321
rect 17865 37312 17877 37315
rect 17828 37284 17877 37312
rect 17828 37272 17834 37284
rect 17865 37281 17877 37284
rect 17911 37281 17923 37315
rect 26329 37315 26387 37321
rect 26329 37312 26341 37315
rect 17865 37275 17923 37281
rect 22020 37284 26341 37312
rect 1581 37247 1639 37253
rect 1581 37213 1593 37247
rect 1627 37244 1639 37247
rect 1762 37244 1768 37256
rect 1627 37216 1768 37244
rect 1627 37213 1639 37216
rect 1581 37207 1639 37213
rect 1762 37204 1768 37216
rect 1820 37204 1826 37256
rect 2498 37244 2504 37256
rect 2459 37216 2504 37244
rect 2498 37204 2504 37216
rect 2556 37204 2562 37256
rect 3234 37244 3240 37256
rect 3195 37216 3240 37244
rect 3234 37204 3240 37216
rect 3292 37204 3298 37256
rect 4341 37247 4399 37253
rect 4341 37213 4353 37247
rect 4387 37244 4399 37247
rect 4706 37244 4712 37256
rect 4387 37216 4712 37244
rect 4387 37213 4399 37216
rect 4341 37207 4399 37213
rect 4706 37204 4712 37216
rect 4764 37204 4770 37256
rect 5077 37247 5135 37253
rect 5077 37213 5089 37247
rect 5123 37213 5135 37247
rect 5810 37244 5816 37256
rect 5771 37216 5816 37244
rect 5077 37207 5135 37213
rect 5092 37176 5120 37207
rect 5810 37204 5816 37216
rect 5868 37204 5874 37256
rect 6917 37247 6975 37253
rect 6917 37213 6929 37247
rect 6963 37244 6975 37247
rect 6963 37216 7328 37244
rect 6963 37213 6975 37216
rect 6917 37207 6975 37213
rect 7006 37176 7012 37188
rect 5092 37148 7012 37176
rect 7006 37136 7012 37148
rect 7064 37136 7070 37188
rect 7300 37176 7328 37216
rect 7374 37204 7380 37256
rect 7432 37244 7438 37256
rect 7653 37247 7711 37253
rect 7653 37244 7665 37247
rect 7432 37216 7665 37244
rect 7432 37204 7438 37216
rect 7653 37213 7665 37216
rect 7699 37213 7711 37247
rect 7653 37207 7711 37213
rect 8389 37247 8447 37253
rect 8389 37213 8401 37247
rect 8435 37244 8447 37247
rect 8570 37244 8576 37256
rect 8435 37216 8576 37244
rect 8435 37213 8447 37216
rect 8389 37207 8447 37213
rect 8570 37204 8576 37216
rect 8628 37204 8634 37256
rect 9493 37247 9551 37253
rect 9493 37213 9505 37247
rect 9539 37244 9551 37247
rect 10229 37247 10287 37253
rect 9539 37216 10180 37244
rect 9539 37213 9551 37216
rect 9493 37207 9551 37213
rect 8294 37176 8300 37188
rect 7300 37148 8300 37176
rect 8294 37136 8300 37148
rect 8352 37136 8358 37188
rect 2314 37108 2320 37120
rect 2275 37080 2320 37108
rect 2314 37068 2320 37080
rect 2372 37068 2378 37120
rect 2866 37068 2872 37120
rect 2924 37108 2930 37120
rect 3053 37111 3111 37117
rect 3053 37108 3065 37111
rect 2924 37080 3065 37108
rect 2924 37068 2930 37080
rect 3053 37077 3065 37080
rect 3099 37077 3111 37111
rect 4154 37108 4160 37120
rect 4115 37080 4160 37108
rect 3053 37071 3111 37077
rect 4154 37068 4160 37080
rect 4212 37068 4218 37120
rect 4893 37111 4951 37117
rect 4893 37077 4905 37111
rect 4939 37108 4951 37111
rect 5074 37108 5080 37120
rect 4939 37080 5080 37108
rect 4939 37077 4951 37080
rect 4893 37071 4951 37077
rect 5074 37068 5080 37080
rect 5132 37068 5138 37120
rect 5626 37108 5632 37120
rect 5587 37080 5632 37108
rect 5626 37068 5632 37080
rect 5684 37068 5690 37120
rect 6730 37108 6736 37120
rect 6691 37080 6736 37108
rect 6730 37068 6736 37080
rect 6788 37068 6794 37120
rect 7282 37068 7288 37120
rect 7340 37108 7346 37120
rect 7469 37111 7527 37117
rect 7469 37108 7481 37111
rect 7340 37080 7481 37108
rect 7340 37068 7346 37080
rect 7469 37077 7481 37080
rect 7515 37077 7527 37111
rect 7469 37071 7527 37077
rect 8205 37111 8263 37117
rect 8205 37077 8217 37111
rect 8251 37108 8263 37111
rect 8386 37108 8392 37120
rect 8251 37080 8392 37108
rect 8251 37077 8263 37080
rect 8205 37071 8263 37077
rect 8386 37068 8392 37080
rect 8444 37068 8450 37120
rect 9309 37111 9367 37117
rect 9309 37077 9321 37111
rect 9355 37108 9367 37111
rect 9490 37108 9496 37120
rect 9355 37080 9496 37108
rect 9355 37077 9367 37080
rect 9309 37071 9367 37077
rect 9490 37068 9496 37080
rect 9548 37068 9554 37120
rect 10042 37108 10048 37120
rect 10003 37080 10048 37108
rect 10042 37068 10048 37080
rect 10100 37068 10106 37120
rect 10152 37108 10180 37216
rect 10229 37213 10241 37247
rect 10275 37213 10287 37247
rect 10229 37207 10287 37213
rect 10244 37176 10272 37207
rect 10318 37204 10324 37256
rect 10376 37244 10382 37256
rect 10689 37247 10747 37253
rect 10689 37244 10701 37247
rect 10376 37216 10701 37244
rect 10376 37204 10382 37216
rect 10689 37213 10701 37216
rect 10735 37213 10747 37247
rect 12066 37244 12072 37256
rect 12027 37216 12072 37244
rect 10689 37207 10747 37213
rect 12066 37204 12072 37216
rect 12124 37204 12130 37256
rect 12526 37244 12532 37256
rect 12487 37216 12532 37244
rect 12526 37204 12532 37216
rect 12584 37204 12590 37256
rect 13538 37244 13544 37256
rect 13499 37216 13544 37244
rect 13538 37204 13544 37216
rect 13596 37204 13602 37256
rect 14642 37244 14648 37256
rect 14603 37216 14648 37244
rect 14642 37204 14648 37216
rect 14700 37204 14706 37256
rect 15378 37244 15384 37256
rect 15339 37216 15384 37244
rect 15378 37204 15384 37216
rect 15436 37204 15442 37256
rect 15838 37244 15844 37256
rect 15799 37216 15844 37244
rect 15838 37204 15844 37216
rect 15896 37204 15902 37256
rect 17405 37247 17463 37253
rect 17405 37213 17417 37247
rect 17451 37244 17463 37247
rect 17678 37244 17684 37256
rect 17451 37216 17684 37244
rect 17451 37213 17463 37216
rect 17405 37207 17463 37213
rect 17678 37204 17684 37216
rect 17736 37204 17742 37256
rect 18141 37247 18199 37253
rect 18141 37213 18153 37247
rect 18187 37213 18199 37247
rect 18141 37207 18199 37213
rect 10410 37176 10416 37188
rect 10244 37148 10416 37176
rect 10410 37136 10416 37148
rect 10468 37136 10474 37188
rect 11054 37176 11060 37188
rect 10520 37148 11060 37176
rect 10520 37108 10548 37148
rect 11054 37136 11060 37148
rect 11112 37136 11118 37188
rect 16850 37136 16856 37188
rect 16908 37176 16914 37188
rect 18156 37176 18184 37207
rect 19334 37204 19340 37256
rect 19392 37244 19398 37256
rect 19613 37247 19671 37253
rect 19613 37244 19625 37247
rect 19392 37216 19625 37244
rect 19392 37204 19398 37216
rect 19613 37213 19625 37216
rect 19659 37244 19671 37247
rect 19978 37244 19984 37256
rect 19659 37216 19984 37244
rect 19659 37213 19671 37216
rect 19613 37207 19671 37213
rect 19978 37204 19984 37216
rect 20036 37204 20042 37256
rect 20162 37204 20168 37256
rect 20220 37244 20226 37256
rect 20257 37247 20315 37253
rect 20257 37244 20269 37247
rect 20220 37216 20269 37244
rect 20220 37204 20226 37216
rect 20257 37213 20269 37216
rect 20303 37213 20315 37247
rect 20257 37207 20315 37213
rect 20438 37204 20444 37256
rect 20496 37244 20502 37256
rect 21085 37247 21143 37253
rect 21085 37244 21097 37247
rect 20496 37216 21097 37244
rect 20496 37204 20502 37216
rect 21085 37213 21097 37216
rect 21131 37213 21143 37247
rect 21085 37207 21143 37213
rect 21174 37204 21180 37256
rect 21232 37244 21238 37256
rect 22020 37253 22048 37284
rect 26329 37281 26341 37284
rect 26375 37281 26387 37315
rect 26329 37275 26387 37281
rect 34238 37272 34244 37324
rect 34296 37312 34302 37324
rect 34701 37315 34759 37321
rect 34701 37312 34713 37315
rect 34296 37284 34713 37312
rect 34296 37272 34302 37284
rect 34701 37281 34713 37284
rect 34747 37281 34759 37315
rect 34701 37275 34759 37281
rect 22005 37247 22063 37253
rect 22005 37244 22017 37247
rect 21232 37216 22017 37244
rect 21232 37204 21238 37216
rect 22005 37213 22017 37216
rect 22051 37213 22063 37247
rect 22005 37207 22063 37213
rect 22094 37204 22100 37256
rect 22152 37244 22158 37256
rect 22649 37247 22707 37253
rect 22649 37244 22661 37247
rect 22152 37216 22661 37244
rect 22152 37204 22158 37216
rect 22649 37213 22661 37216
rect 22695 37213 22707 37247
rect 23290 37244 23296 37256
rect 22649 37207 22707 37213
rect 22940 37216 23296 37244
rect 16908 37148 18184 37176
rect 16908 37136 16914 37148
rect 20806 37136 20812 37188
rect 20864 37176 20870 37188
rect 20864 37148 22094 37176
rect 20864 37136 20870 37148
rect 10152 37080 10548 37108
rect 10873 37111 10931 37117
rect 10873 37077 10885 37111
rect 10919 37108 10931 37111
rect 11146 37108 11152 37120
rect 10919 37080 11152 37108
rect 10919 37077 10931 37080
rect 10873 37071 10931 37077
rect 11146 37068 11152 37080
rect 11204 37068 11210 37120
rect 11698 37068 11704 37120
rect 11756 37108 11762 37120
rect 11885 37111 11943 37117
rect 11885 37108 11897 37111
rect 11756 37080 11897 37108
rect 11756 37068 11762 37080
rect 11885 37077 11897 37080
rect 11931 37077 11943 37111
rect 11885 37071 11943 37077
rect 12713 37111 12771 37117
rect 12713 37077 12725 37111
rect 12759 37108 12771 37111
rect 12802 37108 12808 37120
rect 12759 37080 12808 37108
rect 12759 37077 12771 37080
rect 12713 37071 12771 37077
rect 12802 37068 12808 37080
rect 12860 37068 12866 37120
rect 13354 37108 13360 37120
rect 13315 37080 13360 37108
rect 13354 37068 13360 37080
rect 13412 37068 13418 37120
rect 14458 37108 14464 37120
rect 14419 37080 14464 37108
rect 14458 37068 14464 37080
rect 14516 37068 14522 37120
rect 15194 37108 15200 37120
rect 15155 37080 15200 37108
rect 15194 37068 15200 37080
rect 15252 37068 15258 37120
rect 16025 37111 16083 37117
rect 16025 37077 16037 37111
rect 16071 37108 16083 37111
rect 16114 37108 16120 37120
rect 16071 37080 16120 37108
rect 16071 37077 16083 37080
rect 16025 37071 16083 37077
rect 16114 37068 16120 37080
rect 16172 37068 16178 37120
rect 17218 37108 17224 37120
rect 17179 37080 17224 37108
rect 17218 37068 17224 37080
rect 17276 37068 17282 37120
rect 19797 37111 19855 37117
rect 19797 37077 19809 37111
rect 19843 37108 19855 37111
rect 20346 37108 20352 37120
rect 19843 37080 20352 37108
rect 19843 37077 19855 37080
rect 19797 37071 19855 37077
rect 20346 37068 20352 37080
rect 20404 37068 20410 37120
rect 20898 37108 20904 37120
rect 20859 37080 20904 37108
rect 20898 37068 20904 37080
rect 20956 37068 20962 37120
rect 20990 37068 20996 37120
rect 21048 37108 21054 37120
rect 21821 37111 21879 37117
rect 21821 37108 21833 37111
rect 21048 37080 21833 37108
rect 21048 37068 21054 37080
rect 21821 37077 21833 37080
rect 21867 37077 21879 37111
rect 22066 37108 22094 37148
rect 22186 37136 22192 37188
rect 22244 37176 22250 37188
rect 22940 37176 22968 37216
rect 23290 37204 23296 37216
rect 23348 37204 23354 37256
rect 23658 37204 23664 37256
rect 23716 37244 23722 37256
rect 24397 37247 24455 37253
rect 24397 37244 24409 37247
rect 23716 37216 24409 37244
rect 23716 37204 23722 37216
rect 24397 37213 24409 37216
rect 24443 37213 24455 37247
rect 25130 37244 25136 37256
rect 24397 37207 24455 37213
rect 24504 37216 25136 37244
rect 22244 37148 22968 37176
rect 22244 37136 22250 37148
rect 23382 37136 23388 37188
rect 23440 37176 23446 37188
rect 24504 37176 24532 37216
rect 25130 37204 25136 37216
rect 25188 37204 25194 37256
rect 25225 37247 25283 37253
rect 25225 37213 25237 37247
rect 25271 37213 25283 37247
rect 25225 37207 25283 37213
rect 23440 37148 24532 37176
rect 23440 37136 23446 37148
rect 22465 37111 22523 37117
rect 22465 37108 22477 37111
rect 22066 37080 22477 37108
rect 21821 37071 21879 37077
rect 22465 37077 22477 37080
rect 22511 37077 22523 37111
rect 23106 37108 23112 37120
rect 23067 37080 23112 37108
rect 22465 37071 22523 37077
rect 23106 37068 23112 37080
rect 23164 37068 23170 37120
rect 24581 37111 24639 37117
rect 24581 37077 24593 37111
rect 24627 37108 24639 37111
rect 24670 37108 24676 37120
rect 24627 37080 24676 37108
rect 24627 37077 24639 37080
rect 24581 37071 24639 37077
rect 24670 37068 24676 37080
rect 24728 37068 24734 37120
rect 25038 37108 25044 37120
rect 24999 37080 25044 37108
rect 25038 37068 25044 37080
rect 25096 37068 25102 37120
rect 25130 37068 25136 37120
rect 25188 37108 25194 37120
rect 25240 37108 25268 37207
rect 25314 37204 25320 37256
rect 25372 37244 25378 37256
rect 25869 37247 25927 37253
rect 25869 37244 25881 37247
rect 25372 37216 25881 37244
rect 25372 37204 25378 37216
rect 25869 37213 25881 37216
rect 25915 37244 25927 37247
rect 27430 37244 27436 37256
rect 25915 37216 27436 37244
rect 25915 37213 25927 37216
rect 25869 37207 25927 37213
rect 27430 37204 27436 37216
rect 27488 37204 27494 37256
rect 27525 37247 27583 37253
rect 27525 37213 27537 37247
rect 27571 37244 27583 37247
rect 28074 37244 28080 37256
rect 27571 37216 28080 37244
rect 27571 37213 27583 37216
rect 27525 37207 27583 37213
rect 28074 37204 28080 37216
rect 28132 37204 28138 37256
rect 28261 37247 28319 37253
rect 28261 37213 28273 37247
rect 28307 37213 28319 37247
rect 28261 37207 28319 37213
rect 28997 37247 29055 37253
rect 28997 37213 29009 37247
rect 29043 37244 29055 37247
rect 29270 37244 29276 37256
rect 29043 37216 29276 37244
rect 29043 37213 29055 37216
rect 28997 37207 29055 37213
rect 28276 37176 28304 37207
rect 29270 37204 29276 37216
rect 29328 37204 29334 37256
rect 29825 37247 29883 37253
rect 29825 37213 29837 37247
rect 29871 37244 29883 37247
rect 30374 37244 30380 37256
rect 29871 37216 30380 37244
rect 29871 37213 29883 37216
rect 29825 37207 29883 37213
rect 30374 37204 30380 37216
rect 30432 37204 30438 37256
rect 30561 37247 30619 37253
rect 30561 37213 30573 37247
rect 30607 37244 30619 37247
rect 31110 37244 31116 37256
rect 30607 37216 31116 37244
rect 30607 37213 30619 37216
rect 30561 37207 30619 37213
rect 31110 37204 31116 37216
rect 31168 37204 31174 37256
rect 31297 37247 31355 37253
rect 31297 37213 31309 37247
rect 31343 37244 31355 37247
rect 32214 37244 32220 37256
rect 31343 37216 32220 37244
rect 31343 37213 31355 37216
rect 31297 37207 31355 37213
rect 32214 37204 32220 37216
rect 32272 37204 32278 37256
rect 32398 37244 32404 37256
rect 32359 37216 32404 37244
rect 32398 37204 32404 37216
rect 32456 37204 32462 37256
rect 32490 37204 32496 37256
rect 32548 37244 32554 37256
rect 33137 37247 33195 37253
rect 32548 37216 33088 37244
rect 32548 37204 32554 37216
rect 30098 37176 30104 37188
rect 28276 37148 30104 37176
rect 30098 37136 30104 37148
rect 30156 37136 30162 37188
rect 31570 37136 31576 37188
rect 31628 37176 31634 37188
rect 33060 37176 33088 37216
rect 33137 37213 33149 37247
rect 33183 37244 33195 37247
rect 33873 37247 33931 37253
rect 33183 37216 33824 37244
rect 33183 37213 33195 37216
rect 33137 37207 33195 37213
rect 33796 37176 33824 37216
rect 33873 37213 33885 37247
rect 33919 37244 33931 37247
rect 34974 37244 34980 37256
rect 33919 37216 34980 37244
rect 33919 37213 33931 37216
rect 33873 37207 33931 37213
rect 34974 37204 34980 37216
rect 35032 37204 35038 37256
rect 35345 37247 35403 37253
rect 35345 37213 35357 37247
rect 35391 37244 35403 37247
rect 36078 37244 36084 37256
rect 35391 37216 36084 37244
rect 35391 37213 35403 37216
rect 35345 37207 35403 37213
rect 36078 37204 36084 37216
rect 36136 37204 36142 37256
rect 37553 37247 37611 37253
rect 37553 37213 37565 37247
rect 37599 37244 37611 37247
rect 37599 37216 38148 37244
rect 37599 37213 37611 37216
rect 37553 37207 37611 37213
rect 34790 37176 34796 37188
rect 31628 37148 32996 37176
rect 33060 37148 33732 37176
rect 33796 37148 34796 37176
rect 31628 37136 31634 37148
rect 25188 37080 25268 37108
rect 25188 37068 25194 37080
rect 25314 37068 25320 37120
rect 25372 37108 25378 37120
rect 25685 37111 25743 37117
rect 25685 37108 25697 37111
rect 25372 37080 25697 37108
rect 25372 37068 25378 37080
rect 25685 37077 25697 37080
rect 25731 37077 25743 37111
rect 25685 37071 25743 37077
rect 27154 37068 27160 37120
rect 27212 37108 27218 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 27212 37080 27353 37108
rect 27212 37068 27218 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27341 37071 27399 37077
rect 27706 37068 27712 37120
rect 27764 37108 27770 37120
rect 28077 37111 28135 37117
rect 28077 37108 28089 37111
rect 27764 37080 28089 37108
rect 27764 37068 27770 37080
rect 28077 37077 28089 37080
rect 28123 37077 28135 37111
rect 28077 37071 28135 37077
rect 28258 37068 28264 37120
rect 28316 37108 28322 37120
rect 28813 37111 28871 37117
rect 28813 37108 28825 37111
rect 28316 37080 28825 37108
rect 28316 37068 28322 37080
rect 28813 37077 28825 37080
rect 28859 37077 28871 37111
rect 28813 37071 28871 37077
rect 28994 37068 29000 37120
rect 29052 37108 29058 37120
rect 29641 37111 29699 37117
rect 29641 37108 29653 37111
rect 29052 37080 29653 37108
rect 29052 37068 29058 37080
rect 29641 37077 29653 37080
rect 29687 37077 29699 37111
rect 29641 37071 29699 37077
rect 29914 37068 29920 37120
rect 29972 37108 29978 37120
rect 31113 37111 31171 37117
rect 31113 37108 31125 37111
rect 29972 37080 31125 37108
rect 29972 37068 29978 37080
rect 31113 37077 31125 37080
rect 31159 37077 31171 37111
rect 31113 37071 31171 37077
rect 31386 37068 31392 37120
rect 31444 37108 31450 37120
rect 32968 37117 32996 37148
rect 33704 37117 33732 37148
rect 34790 37136 34796 37148
rect 34848 37136 34854 37188
rect 35618 37185 35624 37188
rect 35612 37139 35624 37185
rect 35676 37176 35682 37188
rect 35676 37148 35712 37176
rect 35866 37148 37412 37176
rect 35618 37136 35624 37139
rect 35676 37136 35682 37148
rect 32217 37111 32275 37117
rect 32217 37108 32229 37111
rect 31444 37080 32229 37108
rect 31444 37068 31450 37080
rect 32217 37077 32229 37080
rect 32263 37077 32275 37111
rect 32217 37071 32275 37077
rect 32953 37111 33011 37117
rect 32953 37077 32965 37111
rect 32999 37077 33011 37111
rect 32953 37071 33011 37077
rect 33689 37111 33747 37117
rect 33689 37077 33701 37111
rect 33735 37077 33747 37111
rect 33689 37071 33747 37077
rect 35342 37068 35348 37120
rect 35400 37108 35406 37120
rect 35866 37108 35894 37148
rect 36722 37108 36728 37120
rect 35400 37080 35894 37108
rect 36683 37080 36728 37108
rect 35400 37068 35406 37080
rect 36722 37068 36728 37080
rect 36780 37068 36786 37120
rect 37384 37117 37412 37148
rect 38120 37117 38148 37216
rect 37369 37111 37427 37117
rect 37369 37077 37381 37111
rect 37415 37077 37427 37111
rect 37369 37071 37427 37077
rect 38105 37111 38163 37117
rect 38105 37077 38117 37111
rect 38151 37108 38163 37111
rect 38286 37108 38292 37120
rect 38151 37080 38292 37108
rect 38151 37077 38163 37080
rect 38105 37071 38163 37077
rect 38286 37068 38292 37080
rect 38344 37068 38350 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1762 36864 1768 36916
rect 1820 36904 1826 36916
rect 1857 36907 1915 36913
rect 1857 36904 1869 36907
rect 1820 36876 1869 36904
rect 1820 36864 1826 36876
rect 1857 36873 1869 36876
rect 1903 36873 1915 36907
rect 1857 36867 1915 36873
rect 2501 36907 2559 36913
rect 2501 36873 2513 36907
rect 2547 36904 2559 36907
rect 3234 36904 3240 36916
rect 2547 36876 3240 36904
rect 2547 36873 2559 36876
rect 2501 36867 2559 36873
rect 3234 36864 3240 36876
rect 3292 36904 3298 36916
rect 3292 36876 4568 36904
rect 3292 36864 3298 36876
rect 3053 36839 3111 36845
rect 3053 36805 3065 36839
rect 3099 36836 3111 36839
rect 3418 36836 3424 36848
rect 3099 36808 3424 36836
rect 3099 36805 3111 36808
rect 3053 36799 3111 36805
rect 3418 36796 3424 36808
rect 3476 36836 3482 36848
rect 3605 36839 3663 36845
rect 3605 36836 3617 36839
rect 3476 36808 3617 36836
rect 3476 36796 3482 36808
rect 3605 36805 3617 36808
rect 3651 36805 3663 36839
rect 4540 36836 4568 36876
rect 4614 36864 4620 36916
rect 4672 36904 4678 36916
rect 4709 36907 4767 36913
rect 4709 36904 4721 36907
rect 4672 36876 4721 36904
rect 4672 36864 4678 36876
rect 4709 36873 4721 36876
rect 4755 36873 4767 36907
rect 4709 36867 4767 36873
rect 6178 36864 6184 36916
rect 6236 36904 6242 36916
rect 6457 36907 6515 36913
rect 6457 36904 6469 36907
rect 6236 36876 6469 36904
rect 6236 36864 6242 36876
rect 6457 36873 6469 36876
rect 6503 36873 6515 36907
rect 6457 36867 6515 36873
rect 7834 36864 7840 36916
rect 7892 36904 7898 36916
rect 8021 36907 8079 36913
rect 8021 36904 8033 36907
rect 7892 36876 8033 36904
rect 7892 36864 7898 36876
rect 8021 36873 8033 36876
rect 8067 36873 8079 36907
rect 8021 36867 8079 36873
rect 8938 36864 8944 36916
rect 8996 36904 9002 36916
rect 9125 36907 9183 36913
rect 9125 36904 9137 36907
rect 8996 36876 9137 36904
rect 8996 36864 9002 36876
rect 9125 36873 9137 36876
rect 9171 36873 9183 36907
rect 9125 36867 9183 36873
rect 10594 36864 10600 36916
rect 10652 36904 10658 36916
rect 10781 36907 10839 36913
rect 10781 36904 10793 36907
rect 10652 36876 10793 36904
rect 10652 36864 10658 36876
rect 10781 36873 10793 36876
rect 10827 36873 10839 36907
rect 12434 36904 12440 36916
rect 12395 36876 12440 36904
rect 10781 36867 10839 36873
rect 12434 36864 12440 36876
rect 12492 36864 12498 36916
rect 13906 36864 13912 36916
rect 13964 36904 13970 36916
rect 14093 36907 14151 36913
rect 14093 36904 14105 36907
rect 13964 36876 14105 36904
rect 13964 36864 13970 36876
rect 14093 36873 14105 36876
rect 14139 36873 14151 36907
rect 14093 36867 14151 36873
rect 15562 36864 15568 36916
rect 15620 36904 15626 36916
rect 15749 36907 15807 36913
rect 15749 36904 15761 36907
rect 15620 36876 15761 36904
rect 15620 36864 15626 36876
rect 15749 36873 15761 36876
rect 15795 36873 15807 36907
rect 15749 36867 15807 36873
rect 16666 36864 16672 36916
rect 16724 36904 16730 36916
rect 16853 36907 16911 36913
rect 16853 36904 16865 36907
rect 16724 36876 16865 36904
rect 16724 36864 16730 36876
rect 16853 36873 16865 36876
rect 16899 36873 16911 36907
rect 16853 36867 16911 36873
rect 19426 36864 19432 36916
rect 19484 36904 19490 36916
rect 19978 36904 19984 36916
rect 19484 36876 19984 36904
rect 19484 36864 19490 36876
rect 19978 36864 19984 36876
rect 20036 36864 20042 36916
rect 20806 36904 20812 36916
rect 20767 36876 20812 36904
rect 20806 36864 20812 36876
rect 20864 36864 20870 36916
rect 20901 36907 20959 36913
rect 20901 36873 20913 36907
rect 20947 36904 20959 36907
rect 21174 36904 21180 36916
rect 20947 36876 21180 36904
rect 20947 36873 20959 36876
rect 20901 36867 20959 36873
rect 21174 36864 21180 36876
rect 21232 36864 21238 36916
rect 21269 36907 21327 36913
rect 21269 36873 21281 36907
rect 21315 36873 21327 36907
rect 23658 36904 23664 36916
rect 23619 36876 23664 36904
rect 21269 36867 21327 36873
rect 9674 36836 9680 36848
rect 4540 36808 9680 36836
rect 3605 36799 3663 36805
rect 9674 36796 9680 36808
rect 9732 36796 9738 36848
rect 13541 36839 13599 36845
rect 13541 36805 13553 36839
rect 13587 36836 13599 36839
rect 14642 36836 14648 36848
rect 13587 36808 14648 36836
rect 13587 36805 13599 36808
rect 13541 36799 13599 36805
rect 14642 36796 14648 36808
rect 14700 36836 14706 36848
rect 18598 36836 18604 36848
rect 14700 36808 18604 36836
rect 14700 36796 14706 36808
rect 18598 36796 18604 36808
rect 18656 36796 18662 36848
rect 19245 36839 19303 36845
rect 19245 36805 19257 36839
rect 19291 36836 19303 36839
rect 20990 36836 20996 36848
rect 19291 36808 20996 36836
rect 19291 36805 19303 36808
rect 19245 36799 19303 36805
rect 20990 36796 20996 36808
rect 21048 36796 21054 36848
rect 4893 36771 4951 36777
rect 4893 36737 4905 36771
rect 4939 36768 4951 36771
rect 5074 36768 5080 36780
rect 4939 36740 5080 36768
rect 4939 36737 4951 36740
rect 4893 36731 4951 36737
rect 5074 36728 5080 36740
rect 5132 36728 5138 36780
rect 6638 36768 6644 36780
rect 6599 36740 6644 36768
rect 6638 36728 6644 36740
rect 6696 36728 6702 36780
rect 8202 36768 8208 36780
rect 8163 36740 8208 36768
rect 8202 36728 8208 36740
rect 8260 36728 8266 36780
rect 9306 36768 9312 36780
rect 9267 36740 9312 36768
rect 9306 36728 9312 36740
rect 9364 36728 9370 36780
rect 10962 36768 10968 36780
rect 10923 36740 10968 36768
rect 10962 36728 10968 36740
rect 11020 36728 11026 36780
rect 12618 36768 12624 36780
rect 12579 36740 12624 36768
rect 12618 36728 12624 36740
rect 12676 36728 12682 36780
rect 14274 36768 14280 36780
rect 14235 36740 14280 36768
rect 14274 36728 14280 36740
rect 14332 36728 14338 36780
rect 15197 36771 15255 36777
rect 15197 36737 15209 36771
rect 15243 36768 15255 36771
rect 15933 36771 15991 36777
rect 15933 36768 15945 36771
rect 15243 36740 15945 36768
rect 15243 36737 15255 36740
rect 15197 36731 15255 36737
rect 15933 36737 15945 36740
rect 15979 36768 15991 36771
rect 16022 36768 16028 36780
rect 15979 36740 16028 36768
rect 15979 36737 15991 36740
rect 15933 36731 15991 36737
rect 16022 36728 16028 36740
rect 16080 36728 16086 36780
rect 17034 36768 17040 36780
rect 16995 36740 17040 36768
rect 17034 36728 17040 36740
rect 17092 36728 17098 36780
rect 17497 36771 17555 36777
rect 17497 36737 17509 36771
rect 17543 36768 17555 36771
rect 17862 36768 17868 36780
rect 17543 36740 17868 36768
rect 17543 36737 17555 36740
rect 17497 36731 17555 36737
rect 17862 36728 17868 36740
rect 17920 36728 17926 36780
rect 18141 36771 18199 36777
rect 18141 36737 18153 36771
rect 18187 36768 18199 36771
rect 19153 36771 19211 36777
rect 18187 36740 18828 36768
rect 18187 36737 18199 36740
rect 18141 36731 18199 36737
rect 3789 36635 3847 36641
rect 3789 36601 3801 36635
rect 3835 36632 3847 36635
rect 6822 36632 6828 36644
rect 3835 36604 6828 36632
rect 3835 36601 3847 36604
rect 3789 36595 3847 36601
rect 6822 36592 6828 36604
rect 6880 36592 6886 36644
rect 18800 36641 18828 36740
rect 19153 36737 19165 36771
rect 19199 36737 19211 36771
rect 21284 36768 21312 36867
rect 23658 36864 23664 36876
rect 23716 36864 23722 36916
rect 24121 36907 24179 36913
rect 24121 36873 24133 36907
rect 24167 36873 24179 36907
rect 24121 36867 24179 36873
rect 24136 36836 24164 36867
rect 25406 36864 25412 36916
rect 25464 36904 25470 36916
rect 25464 36876 26280 36904
rect 25464 36864 25470 36876
rect 22066 36808 24164 36836
rect 21821 36771 21879 36777
rect 21821 36768 21833 36771
rect 21284 36740 21833 36768
rect 19153 36731 19211 36737
rect 21821 36737 21833 36740
rect 21867 36737 21879 36771
rect 22066 36768 22094 36808
rect 24210 36796 24216 36848
rect 24268 36836 24274 36848
rect 24762 36836 24768 36848
rect 24268 36808 24768 36836
rect 24268 36796 24274 36808
rect 24762 36796 24768 36808
rect 24820 36836 24826 36848
rect 26252 36836 26280 36876
rect 28166 36864 28172 36916
rect 28224 36904 28230 36916
rect 28224 36876 30052 36904
rect 28224 36864 28230 36876
rect 29926 36839 29984 36845
rect 29926 36836 29938 36839
rect 24820 36808 25452 36836
rect 26252 36808 29938 36836
rect 24820 36796 24826 36808
rect 21821 36731 21879 36737
rect 21928 36740 22094 36768
rect 23293 36771 23351 36777
rect 18785 36635 18843 36641
rect 18785 36601 18797 36635
rect 18831 36601 18843 36635
rect 19168 36632 19196 36731
rect 19426 36700 19432 36712
rect 19339 36672 19432 36700
rect 19426 36660 19432 36672
rect 19484 36700 19490 36712
rect 20717 36703 20775 36709
rect 20717 36700 20729 36703
rect 19484 36672 20729 36700
rect 19484 36660 19490 36672
rect 20717 36669 20729 36672
rect 20763 36700 20775 36703
rect 21542 36700 21548 36712
rect 20763 36672 21548 36700
rect 20763 36669 20775 36672
rect 20717 36663 20775 36669
rect 21542 36660 21548 36672
rect 21600 36660 21606 36712
rect 20254 36632 20260 36644
rect 19168 36604 20260 36632
rect 18785 36595 18843 36601
rect 20254 36592 20260 36604
rect 20312 36632 20318 36644
rect 21928 36632 21956 36740
rect 23293 36737 23305 36771
rect 23339 36768 23351 36771
rect 23382 36768 23388 36780
rect 23339 36740 23388 36768
rect 23339 36737 23351 36740
rect 23293 36731 23351 36737
rect 23382 36728 23388 36740
rect 23440 36728 23446 36780
rect 25234 36771 25292 36777
rect 25234 36768 25246 36771
rect 23676 36740 25246 36768
rect 23014 36700 23020 36712
rect 22975 36672 23020 36700
rect 23014 36660 23020 36672
rect 23072 36660 23078 36712
rect 23201 36703 23259 36709
rect 23201 36669 23213 36703
rect 23247 36700 23259 36703
rect 23474 36700 23480 36712
rect 23247 36672 23480 36700
rect 23247 36669 23259 36672
rect 23201 36663 23259 36669
rect 23474 36660 23480 36672
rect 23532 36660 23538 36712
rect 20312 36604 21956 36632
rect 22005 36635 22063 36641
rect 20312 36592 20318 36604
rect 22005 36601 22017 36635
rect 22051 36632 22063 36635
rect 23382 36632 23388 36644
rect 22051 36604 23388 36632
rect 22051 36601 22063 36604
rect 22005 36595 22063 36601
rect 23382 36592 23388 36604
rect 23440 36592 23446 36644
rect 5810 36564 5816 36576
rect 5771 36536 5816 36564
rect 5810 36524 5816 36536
rect 5868 36524 5874 36576
rect 7374 36564 7380 36576
rect 7335 36536 7380 36564
rect 7374 36524 7380 36536
rect 7432 36524 7438 36576
rect 10226 36564 10232 36576
rect 10187 36536 10232 36564
rect 10226 36524 10232 36536
rect 10284 36524 10290 36576
rect 11885 36567 11943 36573
rect 11885 36533 11897 36567
rect 11931 36564 11943 36567
rect 12526 36564 12532 36576
rect 11931 36536 12532 36564
rect 11931 36533 11943 36536
rect 11885 36527 11943 36533
rect 12526 36524 12532 36536
rect 12584 36524 12590 36576
rect 17681 36567 17739 36573
rect 17681 36533 17693 36567
rect 17727 36564 17739 36567
rect 17862 36564 17868 36576
rect 17727 36536 17868 36564
rect 17727 36533 17739 36536
rect 17681 36527 17739 36533
rect 17862 36524 17868 36536
rect 17920 36524 17926 36576
rect 18325 36567 18383 36573
rect 18325 36533 18337 36567
rect 18371 36564 18383 36567
rect 23676 36564 23704 36740
rect 25234 36737 25246 36740
rect 25280 36737 25292 36771
rect 25424 36768 25452 36808
rect 29926 36805 29938 36808
rect 29972 36805 29984 36839
rect 30024 36836 30052 36876
rect 30466 36864 30472 36916
rect 30524 36904 30530 36916
rect 30745 36907 30803 36913
rect 30745 36904 30757 36907
rect 30524 36876 30757 36904
rect 30524 36864 30530 36876
rect 30745 36873 30757 36876
rect 30791 36873 30803 36907
rect 30745 36867 30803 36873
rect 34514 36864 34520 36916
rect 34572 36904 34578 36916
rect 35897 36907 35955 36913
rect 35897 36904 35909 36907
rect 34572 36876 35909 36904
rect 34572 36864 34578 36876
rect 35897 36873 35909 36876
rect 35943 36873 35955 36907
rect 35897 36867 35955 36873
rect 37369 36907 37427 36913
rect 37369 36873 37381 36907
rect 37415 36873 37427 36907
rect 37369 36867 37427 36873
rect 33238 36839 33296 36845
rect 33238 36836 33250 36839
rect 30024 36808 33250 36836
rect 29926 36799 29984 36805
rect 33238 36805 33250 36808
rect 33284 36805 33296 36839
rect 33238 36799 33296 36805
rect 35066 36796 35072 36848
rect 35124 36845 35130 36848
rect 35124 36836 35136 36845
rect 37384 36836 37412 36867
rect 35124 36808 35169 36836
rect 35912 36808 37412 36836
rect 35124 36799 35136 36808
rect 35124 36796 35130 36799
rect 35912 36780 35940 36808
rect 26145 36771 26203 36777
rect 26145 36768 26157 36771
rect 25424 36740 26157 36768
rect 25234 36731 25292 36737
rect 26145 36737 26157 36740
rect 26191 36737 26203 36771
rect 28086 36771 28144 36777
rect 28086 36768 28098 36771
rect 26145 36731 26203 36737
rect 26252 36740 28098 36768
rect 25498 36700 25504 36712
rect 25459 36672 25504 36700
rect 25498 36660 25504 36672
rect 25556 36660 25562 36712
rect 26252 36632 26280 36740
rect 28086 36737 28098 36740
rect 28132 36737 28144 36771
rect 30929 36771 30987 36777
rect 28086 36731 28144 36737
rect 29104 36740 30328 36768
rect 28353 36703 28411 36709
rect 28353 36669 28365 36703
rect 28399 36700 28411 36703
rect 28994 36700 29000 36712
rect 28399 36672 29000 36700
rect 28399 36669 28411 36672
rect 28353 36663 28411 36669
rect 28994 36660 29000 36672
rect 29052 36660 29058 36712
rect 25516 36604 26280 36632
rect 18371 36536 23704 36564
rect 18371 36533 18383 36536
rect 18325 36527 18383 36533
rect 23750 36524 23756 36576
rect 23808 36564 23814 36576
rect 25516 36564 25544 36604
rect 26326 36592 26332 36644
rect 26384 36632 26390 36644
rect 26384 36604 27108 36632
rect 26384 36592 26390 36604
rect 25958 36564 25964 36576
rect 23808 36536 25544 36564
rect 25919 36536 25964 36564
rect 23808 36524 23814 36536
rect 25958 36524 25964 36536
rect 26016 36524 26022 36576
rect 26970 36564 26976 36576
rect 26931 36536 26976 36564
rect 26970 36524 26976 36536
rect 27028 36524 27034 36576
rect 27080 36564 27108 36604
rect 28442 36592 28448 36644
rect 28500 36632 28506 36644
rect 28813 36635 28871 36641
rect 28813 36632 28825 36635
rect 28500 36604 28825 36632
rect 28500 36592 28506 36604
rect 28813 36601 28825 36604
rect 28859 36601 28871 36635
rect 28813 36595 28871 36601
rect 29104 36564 29132 36740
rect 30190 36700 30196 36712
rect 30151 36672 30196 36700
rect 30190 36660 30196 36672
rect 30248 36660 30254 36712
rect 30300 36700 30328 36740
rect 30929 36737 30941 36771
rect 30975 36768 30987 36771
rect 31294 36768 31300 36780
rect 30975 36740 31300 36768
rect 30975 36737 30987 36740
rect 30929 36731 30987 36737
rect 31294 36728 31300 36740
rect 31352 36728 31358 36780
rect 35894 36728 35900 36780
rect 35952 36728 35958 36780
rect 36081 36771 36139 36777
rect 36081 36737 36093 36771
rect 36127 36768 36139 36771
rect 36446 36768 36452 36780
rect 36127 36740 36452 36768
rect 36127 36737 36139 36740
rect 36081 36731 36139 36737
rect 36446 36728 36452 36740
rect 36504 36728 36510 36780
rect 37553 36771 37611 36777
rect 37553 36737 37565 36771
rect 37599 36768 37611 36771
rect 38102 36768 38108 36780
rect 37599 36740 38108 36768
rect 37599 36737 37611 36740
rect 37553 36731 37611 36737
rect 38102 36728 38108 36740
rect 38160 36728 38166 36780
rect 33505 36703 33563 36709
rect 30300 36672 31754 36700
rect 31726 36632 31754 36672
rect 33505 36669 33517 36703
rect 33551 36700 33563 36703
rect 33778 36700 33784 36712
rect 33551 36672 33784 36700
rect 33551 36669 33563 36672
rect 33505 36663 33563 36669
rect 33778 36660 33784 36672
rect 33836 36660 33842 36712
rect 35345 36703 35403 36709
rect 35345 36669 35357 36703
rect 35391 36700 35403 36703
rect 35391 36672 36124 36700
rect 35391 36669 35403 36672
rect 35345 36663 35403 36669
rect 36096 36644 36124 36672
rect 32125 36635 32183 36641
rect 32125 36632 32137 36635
rect 31726 36604 32137 36632
rect 32125 36601 32137 36604
rect 32171 36601 32183 36635
rect 32125 36595 32183 36601
rect 35434 36592 35440 36644
rect 35492 36632 35498 36644
rect 35894 36632 35900 36644
rect 35492 36604 35900 36632
rect 35492 36592 35498 36604
rect 35894 36592 35900 36604
rect 35952 36592 35958 36644
rect 36078 36592 36084 36644
rect 36136 36592 36142 36644
rect 27080 36536 29132 36564
rect 29270 36524 29276 36576
rect 29328 36564 29334 36576
rect 31389 36567 31447 36573
rect 31389 36564 31401 36567
rect 29328 36536 31401 36564
rect 29328 36524 29334 36536
rect 31389 36533 31401 36536
rect 31435 36533 31447 36567
rect 33962 36564 33968 36576
rect 33923 36536 33968 36564
rect 31389 36527 31447 36533
rect 33962 36524 33968 36536
rect 34020 36524 34026 36576
rect 34974 36524 34980 36576
rect 35032 36564 35038 36576
rect 36633 36567 36691 36573
rect 36633 36564 36645 36567
rect 35032 36536 36645 36564
rect 35032 36524 35038 36536
rect 36633 36533 36645 36536
rect 36679 36564 36691 36567
rect 37918 36564 37924 36576
rect 36679 36536 37924 36564
rect 36679 36533 36691 36536
rect 36633 36527 36691 36533
rect 37918 36524 37924 36536
rect 37976 36524 37982 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 14274 36320 14280 36372
rect 14332 36360 14338 36372
rect 14461 36363 14519 36369
rect 14461 36360 14473 36363
rect 14332 36332 14473 36360
rect 14332 36320 14338 36332
rect 14461 36329 14473 36332
rect 14507 36360 14519 36363
rect 16574 36360 16580 36372
rect 14507 36332 16580 36360
rect 14507 36329 14519 36332
rect 14461 36323 14519 36329
rect 16574 36320 16580 36332
rect 16632 36320 16638 36372
rect 16945 36363 17003 36369
rect 16945 36329 16957 36363
rect 16991 36360 17003 36363
rect 17770 36360 17776 36372
rect 16991 36332 17776 36360
rect 16991 36329 17003 36332
rect 16945 36323 17003 36329
rect 17770 36320 17776 36332
rect 17828 36320 17834 36372
rect 19426 36360 19432 36372
rect 19387 36332 19432 36360
rect 19426 36320 19432 36332
rect 19484 36320 19490 36372
rect 20162 36360 20168 36372
rect 20123 36332 20168 36360
rect 20162 36320 20168 36332
rect 20220 36320 20226 36372
rect 22741 36363 22799 36369
rect 22741 36329 22753 36363
rect 22787 36360 22799 36363
rect 22787 36332 26740 36360
rect 22787 36329 22799 36332
rect 22741 36323 22799 36329
rect 6638 36252 6644 36304
rect 6696 36292 6702 36304
rect 6825 36295 6883 36301
rect 6825 36292 6837 36295
rect 6696 36264 6837 36292
rect 6696 36252 6702 36264
rect 6825 36261 6837 36264
rect 6871 36292 6883 36295
rect 10042 36292 10048 36304
rect 6871 36264 10048 36292
rect 6871 36261 6883 36264
rect 6825 36255 6883 36261
rect 10042 36252 10048 36264
rect 10100 36252 10106 36304
rect 16393 36295 16451 36301
rect 16393 36261 16405 36295
rect 16439 36292 16451 36295
rect 17678 36292 17684 36304
rect 16439 36264 17684 36292
rect 16439 36261 16451 36264
rect 16393 36255 16451 36261
rect 17678 36252 17684 36264
rect 17736 36252 17742 36304
rect 18693 36295 18751 36301
rect 18693 36261 18705 36295
rect 18739 36292 18751 36295
rect 20070 36292 20076 36304
rect 18739 36264 20076 36292
rect 18739 36261 18751 36264
rect 18693 36255 18751 36261
rect 20070 36252 20076 36264
rect 20128 36252 20134 36304
rect 22097 36295 22155 36301
rect 22097 36261 22109 36295
rect 22143 36292 22155 36295
rect 23385 36295 23443 36301
rect 22143 36264 23244 36292
rect 22143 36261 22155 36264
rect 22097 36255 22155 36261
rect 2498 36184 2504 36236
rect 2556 36224 2562 36236
rect 2685 36227 2743 36233
rect 2685 36224 2697 36227
rect 2556 36196 2697 36224
rect 2556 36184 2562 36196
rect 2685 36193 2697 36196
rect 2731 36224 2743 36227
rect 8754 36224 8760 36236
rect 2731 36196 8760 36224
rect 2731 36193 2743 36196
rect 2685 36187 2743 36193
rect 8754 36184 8760 36196
rect 8812 36184 8818 36236
rect 9306 36184 9312 36236
rect 9364 36224 9370 36236
rect 9493 36227 9551 36233
rect 9493 36224 9505 36227
rect 9364 36196 9505 36224
rect 9364 36184 9370 36196
rect 9493 36193 9505 36196
rect 9539 36224 9551 36227
rect 12710 36224 12716 36236
rect 9539 36196 12716 36224
rect 9539 36193 9551 36196
rect 9493 36187 9551 36193
rect 12710 36184 12716 36196
rect 12768 36184 12774 36236
rect 15289 36227 15347 36233
rect 15289 36193 15301 36227
rect 15335 36224 15347 36227
rect 15378 36224 15384 36236
rect 15335 36196 15384 36224
rect 15335 36193 15347 36196
rect 15289 36187 15347 36193
rect 15378 36184 15384 36196
rect 15436 36224 15442 36236
rect 18414 36224 18420 36236
rect 15436 36196 18420 36224
rect 15436 36184 15442 36196
rect 18414 36184 18420 36196
rect 18472 36184 18478 36236
rect 20622 36224 20628 36236
rect 19352 36196 20628 36224
rect 7377 36159 7435 36165
rect 7377 36125 7389 36159
rect 7423 36156 7435 36159
rect 8294 36156 8300 36168
rect 7423 36128 8300 36156
rect 7423 36125 7435 36128
rect 7377 36119 7435 36125
rect 8294 36116 8300 36128
rect 8352 36156 8358 36168
rect 8938 36156 8944 36168
rect 8352 36128 8944 36156
rect 8352 36116 8358 36128
rect 8938 36116 8944 36128
rect 8996 36116 9002 36168
rect 10410 36156 10416 36168
rect 10323 36128 10416 36156
rect 10410 36116 10416 36128
rect 10468 36156 10474 36168
rect 13170 36156 13176 36168
rect 10468 36128 13176 36156
rect 10468 36116 10474 36128
rect 13170 36116 13176 36128
rect 13228 36116 13234 36168
rect 13538 36156 13544 36168
rect 13451 36128 13544 36156
rect 13538 36116 13544 36128
rect 13596 36156 13602 36168
rect 15746 36156 15752 36168
rect 13596 36128 15752 36156
rect 13596 36116 13602 36128
rect 15746 36116 15752 36128
rect 15804 36116 15810 36168
rect 17497 36159 17555 36165
rect 17497 36125 17509 36159
rect 17543 36156 17555 36159
rect 18509 36159 18567 36165
rect 18509 36156 18521 36159
rect 17543 36128 18521 36156
rect 17543 36125 17555 36128
rect 17497 36119 17555 36125
rect 18509 36125 18521 36128
rect 18555 36156 18567 36159
rect 18874 36156 18880 36168
rect 18555 36128 18880 36156
rect 18555 36125 18567 36128
rect 18509 36119 18567 36125
rect 18874 36116 18880 36128
rect 18932 36116 18938 36168
rect 19352 36165 19380 36196
rect 20622 36184 20628 36196
rect 20680 36224 20686 36236
rect 20717 36227 20775 36233
rect 20717 36224 20729 36227
rect 20680 36196 20729 36224
rect 20680 36184 20686 36196
rect 20717 36193 20729 36196
rect 20763 36193 20775 36227
rect 21542 36224 21548 36236
rect 21503 36196 21548 36224
rect 20717 36187 20775 36193
rect 21542 36184 21548 36196
rect 21600 36184 21606 36236
rect 21637 36227 21695 36233
rect 21637 36193 21649 36227
rect 21683 36224 21695 36227
rect 23106 36224 23112 36236
rect 21683 36196 23112 36224
rect 21683 36193 21695 36196
rect 21637 36187 21695 36193
rect 23106 36184 23112 36196
rect 23164 36184 23170 36236
rect 19337 36159 19395 36165
rect 19337 36125 19349 36159
rect 19383 36125 19395 36159
rect 22370 36156 22376 36168
rect 19337 36119 19395 36125
rect 20640 36128 22376 36156
rect 5629 36091 5687 36097
rect 5629 36057 5641 36091
rect 5675 36088 5687 36091
rect 7006 36088 7012 36100
rect 5675 36060 7012 36088
rect 5675 36057 5687 36060
rect 5629 36051 5687 36057
rect 7006 36048 7012 36060
rect 7064 36088 7070 36100
rect 7558 36088 7564 36100
rect 7064 36060 7564 36088
rect 7064 36048 7070 36060
rect 7558 36048 7564 36060
rect 7616 36048 7622 36100
rect 10962 36048 10968 36100
rect 11020 36088 11026 36100
rect 11149 36091 11207 36097
rect 11149 36088 11161 36091
rect 11020 36060 11161 36088
rect 11020 36048 11026 36060
rect 11149 36057 11161 36060
rect 11195 36088 11207 36091
rect 13630 36088 13636 36100
rect 11195 36060 13636 36088
rect 11195 36057 11207 36060
rect 11149 36051 11207 36057
rect 13630 36048 13636 36060
rect 13688 36048 13694 36100
rect 18049 36091 18107 36097
rect 18049 36057 18061 36091
rect 18095 36088 18107 36091
rect 20438 36088 20444 36100
rect 18095 36060 20444 36088
rect 18095 36057 18107 36060
rect 18049 36051 18107 36057
rect 20438 36048 20444 36060
rect 20496 36048 20502 36100
rect 20640 36097 20668 36128
rect 22370 36116 22376 36128
rect 22428 36116 22434 36168
rect 22554 36156 22560 36168
rect 22515 36128 22560 36156
rect 22554 36116 22560 36128
rect 22612 36116 22618 36168
rect 23216 36165 23244 36264
rect 23385 36261 23397 36295
rect 23431 36292 23443 36295
rect 23750 36292 23756 36304
rect 23431 36264 23756 36292
rect 23431 36261 23443 36264
rect 23385 36255 23443 36261
rect 23750 36252 23756 36264
rect 23808 36252 23814 36304
rect 23474 36184 23480 36236
rect 23532 36224 23538 36236
rect 25314 36224 25320 36236
rect 23532 36196 25320 36224
rect 23532 36184 23538 36196
rect 25314 36184 25320 36196
rect 25372 36184 25378 36236
rect 23201 36159 23259 36165
rect 23201 36125 23213 36159
rect 23247 36125 23259 36159
rect 24394 36156 24400 36168
rect 24355 36128 24400 36156
rect 23201 36119 23259 36125
rect 24394 36116 24400 36128
rect 24452 36116 24458 36168
rect 25498 36116 25504 36168
rect 25556 36156 25562 36168
rect 26513 36159 26571 36165
rect 26513 36156 26525 36159
rect 25556 36128 26525 36156
rect 25556 36116 25562 36128
rect 26513 36125 26525 36128
rect 26559 36125 26571 36159
rect 26712 36156 26740 36332
rect 27430 36320 27436 36372
rect 27488 36360 27494 36372
rect 29549 36363 29607 36369
rect 29549 36360 29561 36363
rect 27488 36332 29561 36360
rect 27488 36320 27494 36332
rect 29549 36329 29561 36332
rect 29595 36329 29607 36363
rect 29549 36323 29607 36329
rect 36538 36320 36544 36372
rect 36596 36360 36602 36372
rect 37185 36363 37243 36369
rect 37185 36360 37197 36363
rect 36596 36332 37197 36360
rect 36596 36320 36602 36332
rect 37185 36329 37197 36332
rect 37231 36329 37243 36363
rect 37185 36323 37243 36329
rect 37090 36252 37096 36304
rect 37148 36292 37154 36304
rect 37921 36295 37979 36301
rect 37921 36292 37933 36295
rect 37148 36264 37933 36292
rect 37148 36252 37154 36264
rect 37921 36261 37933 36264
rect 37967 36261 37979 36295
rect 37921 36255 37979 36261
rect 29454 36184 29460 36236
rect 29512 36224 29518 36236
rect 33778 36224 33784 36236
rect 29512 36196 30328 36224
rect 33739 36196 33784 36224
rect 29512 36184 29518 36196
rect 28546 36159 28604 36165
rect 28546 36156 28558 36159
rect 26712 36128 28558 36156
rect 26513 36119 26571 36125
rect 28546 36125 28558 36128
rect 28592 36125 28604 36159
rect 28546 36119 28604 36125
rect 28813 36159 28871 36165
rect 28813 36125 28825 36159
rect 28859 36156 28871 36159
rect 28994 36156 29000 36168
rect 28859 36128 29000 36156
rect 28859 36125 28871 36128
rect 28813 36119 28871 36125
rect 28994 36116 29000 36128
rect 29052 36156 29058 36168
rect 30006 36156 30012 36168
rect 29052 36128 30012 36156
rect 29052 36116 29058 36128
rect 30006 36116 30012 36128
rect 30064 36156 30070 36168
rect 30190 36156 30196 36168
rect 30064 36128 30196 36156
rect 30064 36116 30070 36128
rect 30190 36116 30196 36128
rect 30248 36116 30254 36168
rect 30300 36156 30328 36196
rect 33778 36184 33784 36196
rect 33836 36184 33842 36236
rect 32398 36156 32404 36168
rect 30300 36128 32404 36156
rect 32398 36116 32404 36128
rect 32456 36156 32462 36168
rect 34238 36156 34244 36168
rect 32456 36128 34244 36156
rect 32456 36116 32462 36128
rect 34238 36116 34244 36128
rect 34296 36116 34302 36168
rect 35161 36159 35219 36165
rect 35161 36125 35173 36159
rect 35207 36156 35219 36159
rect 37001 36159 37059 36165
rect 37001 36156 37013 36159
rect 35207 36128 35894 36156
rect 35207 36125 35219 36128
rect 35161 36119 35219 36125
rect 20625 36091 20683 36097
rect 20625 36057 20637 36091
rect 20671 36057 20683 36091
rect 20625 36051 20683 36057
rect 21266 36048 21272 36100
rect 21324 36088 21330 36100
rect 21726 36088 21732 36100
rect 21324 36060 21732 36088
rect 21324 36048 21330 36060
rect 21726 36048 21732 36060
rect 21784 36048 21790 36100
rect 22094 36048 22100 36100
rect 22152 36088 22158 36100
rect 25958 36088 25964 36100
rect 22152 36060 25964 36088
rect 22152 36048 22158 36060
rect 25958 36048 25964 36060
rect 26016 36048 26022 36100
rect 26234 36088 26240 36100
rect 26292 36097 26298 36100
rect 26204 36060 26240 36088
rect 26234 36048 26240 36060
rect 26292 36051 26304 36097
rect 26292 36048 26298 36051
rect 30282 36048 30288 36100
rect 30340 36088 30346 36100
rect 30438 36091 30496 36097
rect 30438 36088 30450 36091
rect 30340 36060 30450 36088
rect 30340 36048 30346 36060
rect 30438 36057 30450 36060
rect 30484 36057 30496 36091
rect 30438 36051 30496 36057
rect 31846 36048 31852 36100
rect 31904 36088 31910 36100
rect 35434 36097 35440 36100
rect 33514 36091 33572 36097
rect 33514 36088 33526 36091
rect 31904 36060 33526 36088
rect 31904 36048 31910 36060
rect 33514 36057 33526 36060
rect 33560 36057 33572 36091
rect 33514 36051 33572 36057
rect 35428 36051 35440 36097
rect 35492 36088 35498 36100
rect 35866 36088 35894 36128
rect 36556 36128 37013 36156
rect 36078 36088 36084 36100
rect 35492 36060 35528 36088
rect 35866 36060 36084 36088
rect 35434 36048 35440 36051
rect 35492 36048 35498 36060
rect 36078 36048 36084 36060
rect 36136 36048 36142 36100
rect 36556 36032 36584 36128
rect 37001 36125 37013 36128
rect 37047 36125 37059 36159
rect 37734 36156 37740 36168
rect 37695 36128 37740 36156
rect 37001 36119 37059 36125
rect 37734 36116 37740 36128
rect 37792 36116 37798 36168
rect 4525 36023 4583 36029
rect 4525 35989 4537 36023
rect 4571 36020 4583 36023
rect 4706 36020 4712 36032
rect 4571 35992 4712 36020
rect 4571 35989 4583 35992
rect 4525 35983 4583 35989
rect 4706 35980 4712 35992
rect 4764 35980 4770 36032
rect 5074 36020 5080 36032
rect 5035 35992 5080 36020
rect 5074 35980 5080 35992
rect 5132 35980 5138 36032
rect 8202 35980 8208 36032
rect 8260 36020 8266 36032
rect 8389 36023 8447 36029
rect 8389 36020 8401 36023
rect 8260 35992 8401 36020
rect 8260 35980 8266 35992
rect 8389 35989 8401 35992
rect 8435 36020 8447 36023
rect 11422 36020 11428 36032
rect 8435 35992 11428 36020
rect 8435 35989 8447 35992
rect 8389 35983 8447 35989
rect 11422 35980 11428 35992
rect 11480 35980 11486 36032
rect 12066 35980 12072 36032
rect 12124 36020 12130 36032
rect 12161 36023 12219 36029
rect 12161 36020 12173 36023
rect 12124 35992 12173 36020
rect 12124 35980 12130 35992
rect 12161 35989 12173 35992
rect 12207 35989 12219 36023
rect 12161 35983 12219 35989
rect 12618 35980 12624 36032
rect 12676 36020 12682 36032
rect 12805 36023 12863 36029
rect 12805 36020 12817 36023
rect 12676 35992 12817 36020
rect 12676 35980 12682 35992
rect 12805 35989 12817 35992
rect 12851 36020 12863 36023
rect 13262 36020 13268 36032
rect 12851 35992 13268 36020
rect 12851 35989 12863 35992
rect 12805 35983 12863 35989
rect 13262 35980 13268 35992
rect 13320 35980 13326 36032
rect 15838 36020 15844 36032
rect 15751 35992 15844 36020
rect 15838 35980 15844 35992
rect 15896 36020 15902 36032
rect 16298 36020 16304 36032
rect 15896 35992 16304 36020
rect 15896 35980 15902 35992
rect 16298 35980 16304 35992
rect 16356 35980 16362 36032
rect 20533 36023 20591 36029
rect 20533 35989 20545 36023
rect 20579 36020 20591 36023
rect 21082 36020 21088 36032
rect 20579 35992 21088 36020
rect 20579 35989 20591 35992
rect 20533 35983 20591 35989
rect 21082 35980 21088 35992
rect 21140 35980 21146 36032
rect 24578 36020 24584 36032
rect 24539 35992 24584 36020
rect 24578 35980 24584 35992
rect 24636 35980 24642 36032
rect 24854 35980 24860 36032
rect 24912 36020 24918 36032
rect 25133 36023 25191 36029
rect 25133 36020 25145 36023
rect 24912 35992 25145 36020
rect 24912 35980 24918 35992
rect 25133 35989 25145 35992
rect 25179 35989 25191 36023
rect 25133 35983 25191 35989
rect 25222 35980 25228 36032
rect 25280 36020 25286 36032
rect 27433 36023 27491 36029
rect 27433 36020 27445 36023
rect 25280 35992 27445 36020
rect 25280 35980 25286 35992
rect 27433 35989 27445 35992
rect 27479 35989 27491 36023
rect 27433 35983 27491 35989
rect 27706 35980 27712 36032
rect 27764 36020 27770 36032
rect 31573 36023 31631 36029
rect 31573 36020 31585 36023
rect 27764 35992 31585 36020
rect 27764 35980 27770 35992
rect 31573 35989 31585 35992
rect 31619 35989 31631 36023
rect 31573 35983 31631 35989
rect 31662 35980 31668 36032
rect 31720 36020 31726 36032
rect 32401 36023 32459 36029
rect 32401 36020 32413 36023
rect 31720 35992 32413 36020
rect 31720 35980 31726 35992
rect 32401 35989 32413 35992
rect 32447 35989 32459 36023
rect 36538 36020 36544 36032
rect 36499 35992 36544 36020
rect 32401 35983 32459 35989
rect 36538 35980 36544 35992
rect 36596 35980 36602 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 17218 35816 17224 35828
rect 17179 35788 17224 35816
rect 17218 35776 17224 35788
rect 17276 35776 17282 35828
rect 17865 35819 17923 35825
rect 17865 35785 17877 35819
rect 17911 35816 17923 35819
rect 17954 35816 17960 35828
rect 17911 35788 17960 35816
rect 17911 35785 17923 35788
rect 17865 35779 17923 35785
rect 17954 35776 17960 35788
rect 18012 35776 18018 35828
rect 18509 35819 18567 35825
rect 18509 35785 18521 35819
rect 18555 35816 18567 35819
rect 19334 35816 19340 35828
rect 18555 35788 19340 35816
rect 18555 35785 18567 35788
rect 18509 35779 18567 35785
rect 19334 35776 19340 35788
rect 19392 35776 19398 35828
rect 21082 35816 21088 35828
rect 21043 35788 21088 35816
rect 21082 35776 21088 35788
rect 21140 35776 21146 35828
rect 22094 35776 22100 35828
rect 22152 35816 22158 35828
rect 22554 35816 22560 35828
rect 22152 35788 22197 35816
rect 22515 35788 22560 35816
rect 22152 35776 22158 35788
rect 22554 35776 22560 35788
rect 22612 35776 22618 35828
rect 23753 35819 23811 35825
rect 23753 35785 23765 35819
rect 23799 35816 23811 35819
rect 24394 35816 24400 35828
rect 23799 35788 24400 35816
rect 23799 35785 23811 35788
rect 23753 35779 23811 35785
rect 24394 35776 24400 35788
rect 24452 35776 24458 35828
rect 26973 35819 27031 35825
rect 26973 35816 26985 35819
rect 25148 35788 26985 35816
rect 13357 35751 13415 35757
rect 13357 35717 13369 35751
rect 13403 35748 13415 35751
rect 13446 35748 13452 35760
rect 13403 35720 13452 35748
rect 13403 35717 13415 35720
rect 13357 35711 13415 35717
rect 13446 35708 13452 35720
rect 13504 35708 13510 35760
rect 19245 35751 19303 35757
rect 19245 35717 19257 35751
rect 19291 35748 19303 35751
rect 23293 35751 23351 35757
rect 19291 35720 23244 35748
rect 19291 35717 19303 35720
rect 19245 35711 19303 35717
rect 13722 35680 13728 35692
rect 13683 35652 13728 35680
rect 13722 35640 13728 35652
rect 13780 35640 13786 35692
rect 13817 35683 13875 35689
rect 13817 35649 13829 35683
rect 13863 35680 13875 35683
rect 14553 35683 14611 35689
rect 14553 35680 14565 35683
rect 13863 35652 14565 35680
rect 13863 35649 13875 35652
rect 13817 35643 13875 35649
rect 14553 35649 14565 35652
rect 14599 35649 14611 35683
rect 14553 35643 14611 35649
rect 15197 35683 15255 35689
rect 15197 35649 15209 35683
rect 15243 35680 15255 35683
rect 16206 35680 16212 35692
rect 15243 35652 16212 35680
rect 15243 35649 15255 35652
rect 15197 35643 15255 35649
rect 16206 35640 16212 35652
rect 16264 35680 16270 35692
rect 16264 35652 19288 35680
rect 16264 35640 16270 35652
rect 11882 35572 11888 35624
rect 11940 35612 11946 35624
rect 13449 35615 13507 35621
rect 13449 35612 13461 35615
rect 11940 35584 13461 35612
rect 11940 35572 11946 35584
rect 13449 35581 13461 35584
rect 13495 35581 13507 35615
rect 14734 35612 14740 35624
rect 14695 35584 14740 35612
rect 13449 35575 13507 35581
rect 14734 35572 14740 35584
rect 14792 35572 14798 35624
rect 14826 35572 14832 35624
rect 14884 35612 14890 35624
rect 16666 35612 16672 35624
rect 14884 35584 16672 35612
rect 14884 35572 14890 35584
rect 16666 35572 16672 35584
rect 16724 35572 16730 35624
rect 19153 35615 19211 35621
rect 19153 35581 19165 35615
rect 19199 35581 19211 35615
rect 19260 35612 19288 35652
rect 19334 35640 19340 35692
rect 19392 35680 19398 35692
rect 19392 35652 19437 35680
rect 19392 35640 19398 35652
rect 19978 35640 19984 35692
rect 20036 35680 20042 35692
rect 20165 35683 20223 35689
rect 20165 35680 20177 35683
rect 20036 35652 20177 35680
rect 20036 35640 20042 35652
rect 20165 35649 20177 35652
rect 20211 35649 20223 35683
rect 20165 35643 20223 35649
rect 20438 35640 20444 35692
rect 20496 35680 20502 35692
rect 22189 35683 22247 35689
rect 20496 35652 21312 35680
rect 20496 35640 20502 35652
rect 19260 35584 21220 35612
rect 19153 35575 19211 35581
rect 19168 35544 19196 35575
rect 19426 35544 19432 35556
rect 19168 35516 19432 35544
rect 19426 35504 19432 35516
rect 19484 35504 19490 35556
rect 8570 35476 8576 35488
rect 8531 35448 8576 35476
rect 8570 35436 8576 35448
rect 8628 35436 8634 35488
rect 9677 35479 9735 35485
rect 9677 35445 9689 35479
rect 9723 35476 9735 35479
rect 11054 35476 11060 35488
rect 9723 35448 11060 35476
rect 9723 35445 9735 35448
rect 9677 35439 9735 35445
rect 11054 35436 11060 35448
rect 11112 35436 11118 35488
rect 13538 35476 13544 35488
rect 13499 35448 13544 35476
rect 13538 35436 13544 35448
rect 13596 35436 13602 35488
rect 13998 35436 14004 35488
rect 14056 35476 14062 35488
rect 16482 35476 16488 35488
rect 14056 35448 16488 35476
rect 14056 35436 14062 35448
rect 16482 35436 16488 35448
rect 16540 35436 16546 35488
rect 19705 35479 19763 35485
rect 19705 35445 19717 35479
rect 19751 35476 19763 35479
rect 19794 35476 19800 35488
rect 19751 35448 19800 35476
rect 19751 35445 19763 35448
rect 19705 35439 19763 35445
rect 19794 35436 19800 35448
rect 19852 35436 19858 35488
rect 20349 35479 20407 35485
rect 20349 35445 20361 35479
rect 20395 35476 20407 35479
rect 21082 35476 21088 35488
rect 20395 35448 21088 35476
rect 20395 35445 20407 35448
rect 20349 35439 20407 35445
rect 21082 35436 21088 35448
rect 21140 35436 21146 35488
rect 21192 35476 21220 35584
rect 21284 35544 21312 35652
rect 22189 35649 22201 35683
rect 22235 35680 22247 35683
rect 22738 35680 22744 35692
rect 22235 35652 22744 35680
rect 22235 35649 22247 35652
rect 22189 35643 22247 35649
rect 22738 35640 22744 35652
rect 22796 35640 22802 35692
rect 21542 35572 21548 35624
rect 21600 35612 21606 35624
rect 21913 35615 21971 35621
rect 21913 35612 21925 35615
rect 21600 35584 21925 35612
rect 21600 35572 21606 35584
rect 21913 35581 21925 35584
rect 21959 35612 21971 35615
rect 23106 35612 23112 35624
rect 21959 35584 23112 35612
rect 21959 35581 21971 35584
rect 21913 35575 21971 35581
rect 23106 35572 23112 35584
rect 23164 35572 23170 35624
rect 23216 35612 23244 35720
rect 23293 35717 23305 35751
rect 23339 35748 23351 35751
rect 25038 35748 25044 35760
rect 23339 35720 25044 35748
rect 23339 35717 23351 35720
rect 23293 35711 23351 35717
rect 25038 35708 25044 35720
rect 25096 35708 25102 35760
rect 23382 35680 23388 35692
rect 23343 35652 23388 35680
rect 23382 35640 23388 35652
rect 23440 35640 23446 35692
rect 25148 35680 25176 35788
rect 26973 35785 26985 35788
rect 27019 35785 27031 35819
rect 26973 35779 27031 35785
rect 30374 35776 30380 35828
rect 30432 35816 30438 35828
rect 30561 35819 30619 35825
rect 30561 35816 30573 35819
rect 30432 35788 30573 35816
rect 30432 35776 30438 35788
rect 30561 35785 30573 35788
rect 30607 35816 30619 35819
rect 30607 35788 31754 35816
rect 30607 35785 30619 35788
rect 30561 35779 30619 35785
rect 26050 35708 26056 35760
rect 26108 35748 26114 35760
rect 26108 35720 27200 35748
rect 26108 35708 26114 35720
rect 25314 35680 25320 35692
rect 25372 35689 25378 35692
rect 23492 35652 25176 35680
rect 25284 35652 25320 35680
rect 23492 35612 23520 35652
rect 25314 35640 25320 35652
rect 25372 35643 25384 35689
rect 25372 35640 25378 35643
rect 25498 35640 25504 35692
rect 25556 35680 25562 35692
rect 25593 35683 25651 35689
rect 25593 35680 25605 35683
rect 25556 35652 25605 35680
rect 25556 35640 25562 35652
rect 25593 35649 25605 35652
rect 25639 35649 25651 35683
rect 25593 35643 25651 35649
rect 25682 35640 25688 35692
rect 25740 35680 25746 35692
rect 27172 35689 27200 35720
rect 26237 35683 26295 35689
rect 26237 35680 26249 35683
rect 25740 35652 26249 35680
rect 25740 35640 25746 35652
rect 26237 35649 26249 35652
rect 26283 35649 26295 35683
rect 26237 35643 26295 35649
rect 27157 35683 27215 35689
rect 27157 35649 27169 35683
rect 27203 35680 27215 35683
rect 27890 35680 27896 35692
rect 27203 35652 27896 35680
rect 27203 35649 27215 35652
rect 27157 35643 27215 35649
rect 23216 35584 23520 35612
rect 26252 35612 26280 35643
rect 27890 35640 27896 35652
rect 27948 35640 27954 35692
rect 27982 35640 27988 35692
rect 28040 35680 28046 35692
rect 29282 35683 29340 35689
rect 29282 35680 29294 35683
rect 28040 35652 29294 35680
rect 28040 35640 28046 35652
rect 29282 35649 29294 35652
rect 29328 35649 29340 35683
rect 29282 35643 29340 35649
rect 27617 35615 27675 35621
rect 27617 35612 27629 35615
rect 26252 35584 27629 35612
rect 27617 35581 27629 35584
rect 27663 35581 27675 35615
rect 27617 35575 27675 35581
rect 29549 35615 29607 35621
rect 29549 35581 29561 35615
rect 29595 35612 29607 35615
rect 30006 35612 30012 35624
rect 29595 35584 30012 35612
rect 29595 35581 29607 35584
rect 29549 35575 29607 35581
rect 30006 35572 30012 35584
rect 30064 35572 30070 35624
rect 24213 35547 24271 35553
rect 24213 35544 24225 35547
rect 21284 35516 24225 35544
rect 24213 35513 24225 35516
rect 24259 35513 24271 35547
rect 31726 35544 31754 35788
rect 32674 35776 32680 35828
rect 32732 35816 32738 35828
rect 32861 35819 32919 35825
rect 32861 35816 32873 35819
rect 32732 35788 32873 35816
rect 32732 35776 32738 35788
rect 32861 35785 32873 35788
rect 32907 35785 32919 35819
rect 32861 35779 32919 35785
rect 33226 35776 33232 35828
rect 33284 35816 33290 35828
rect 33597 35819 33655 35825
rect 33597 35816 33609 35819
rect 33284 35788 33609 35816
rect 33284 35776 33290 35788
rect 33597 35785 33609 35788
rect 33643 35785 33655 35819
rect 33597 35779 33655 35785
rect 33870 35776 33876 35828
rect 33928 35816 33934 35828
rect 34333 35819 34391 35825
rect 34333 35816 34345 35819
rect 33928 35788 34345 35816
rect 33928 35776 33934 35788
rect 34333 35785 34345 35788
rect 34379 35785 34391 35819
rect 34333 35779 34391 35785
rect 35986 35776 35992 35828
rect 36044 35816 36050 35828
rect 36173 35819 36231 35825
rect 36173 35816 36185 35819
rect 36044 35788 36185 35816
rect 36044 35776 36050 35788
rect 36173 35785 36185 35788
rect 36219 35785 36231 35819
rect 36173 35779 36231 35785
rect 37642 35776 37648 35828
rect 37700 35816 37706 35828
rect 37829 35819 37887 35825
rect 37829 35816 37841 35819
rect 37700 35788 37841 35816
rect 37700 35776 37706 35788
rect 37829 35785 37841 35788
rect 37875 35785 37887 35819
rect 37829 35779 37887 35785
rect 33045 35683 33103 35689
rect 33045 35649 33057 35683
rect 33091 35649 33103 35683
rect 33045 35643 33103 35649
rect 33781 35683 33839 35689
rect 33781 35649 33793 35683
rect 33827 35680 33839 35683
rect 34517 35683 34575 35689
rect 33827 35652 34468 35680
rect 33827 35649 33839 35652
rect 33781 35643 33839 35649
rect 33060 35612 33088 35643
rect 34054 35612 34060 35624
rect 33060 35584 34060 35612
rect 34054 35572 34060 35584
rect 34112 35572 34118 35624
rect 34440 35612 34468 35652
rect 34517 35649 34529 35683
rect 34563 35680 34575 35683
rect 36170 35680 36176 35692
rect 34563 35652 36176 35680
rect 34563 35649 34575 35652
rect 34517 35643 34575 35649
rect 36170 35640 36176 35652
rect 36228 35640 36234 35692
rect 36357 35683 36415 35689
rect 36357 35649 36369 35683
rect 36403 35680 36415 35683
rect 36722 35680 36728 35692
rect 36403 35652 36728 35680
rect 36403 35649 36415 35652
rect 36357 35643 36415 35649
rect 35342 35612 35348 35624
rect 34440 35584 35348 35612
rect 35342 35572 35348 35584
rect 35400 35572 35406 35624
rect 36372 35612 36400 35643
rect 36722 35640 36728 35652
rect 36780 35640 36786 35692
rect 37642 35640 37648 35692
rect 37700 35680 37706 35692
rect 38013 35683 38071 35689
rect 38013 35680 38025 35683
rect 37700 35652 38025 35680
rect 37700 35640 37706 35652
rect 38013 35649 38025 35652
rect 38059 35649 38071 35683
rect 38013 35643 38071 35649
rect 35912 35584 36400 35612
rect 32858 35544 32864 35556
rect 31726 35516 32864 35544
rect 24213 35507 24271 35513
rect 32858 35504 32864 35516
rect 32916 35504 32922 35556
rect 35912 35488 35940 35584
rect 24854 35476 24860 35488
rect 21192 35448 24860 35476
rect 24854 35436 24860 35448
rect 24912 35436 24918 35488
rect 26050 35476 26056 35488
rect 26011 35448 26056 35476
rect 26050 35436 26056 35448
rect 26108 35436 26114 35488
rect 27614 35436 27620 35488
rect 27672 35476 27678 35488
rect 28169 35479 28227 35485
rect 28169 35476 28181 35479
rect 27672 35448 28181 35476
rect 27672 35436 27678 35448
rect 28169 35445 28181 35448
rect 28215 35445 28227 35479
rect 30098 35476 30104 35488
rect 30059 35448 30104 35476
rect 28169 35439 28227 35445
rect 30098 35436 30104 35448
rect 30156 35436 30162 35488
rect 31110 35476 31116 35488
rect 31071 35448 31116 35476
rect 31110 35436 31116 35448
rect 31168 35436 31174 35488
rect 32122 35476 32128 35488
rect 32083 35448 32128 35476
rect 32122 35436 32128 35448
rect 32180 35436 32186 35488
rect 34698 35436 34704 35488
rect 34756 35476 34762 35488
rect 34977 35479 35035 35485
rect 34977 35476 34989 35479
rect 34756 35448 34989 35476
rect 34756 35436 34762 35448
rect 34977 35445 34989 35448
rect 35023 35445 35035 35479
rect 34977 35439 35035 35445
rect 35621 35479 35679 35485
rect 35621 35445 35633 35479
rect 35667 35476 35679 35479
rect 35894 35476 35900 35488
rect 35667 35448 35900 35476
rect 35667 35445 35679 35448
rect 35621 35439 35679 35445
rect 35894 35436 35900 35448
rect 35952 35436 35958 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 10870 35232 10876 35284
rect 10928 35272 10934 35284
rect 10928 35244 14596 35272
rect 10928 35232 10934 35244
rect 13814 35164 13820 35216
rect 13872 35204 13878 35216
rect 14461 35207 14519 35213
rect 14461 35204 14473 35207
rect 13872 35176 14473 35204
rect 13872 35164 13878 35176
rect 14461 35173 14473 35176
rect 14507 35173 14519 35207
rect 14568 35204 14596 35244
rect 14734 35232 14740 35284
rect 14792 35272 14798 35284
rect 15381 35275 15439 35281
rect 15381 35272 15393 35275
rect 14792 35244 15393 35272
rect 14792 35232 14798 35244
rect 15381 35241 15393 35244
rect 15427 35241 15439 35275
rect 19334 35272 19340 35284
rect 15381 35235 15439 35241
rect 16132 35244 16436 35272
rect 19295 35244 19340 35272
rect 15654 35204 15660 35216
rect 14568 35176 15660 35204
rect 14461 35167 14519 35173
rect 15654 35164 15660 35176
rect 15712 35164 15718 35216
rect 12894 35096 12900 35148
rect 12952 35136 12958 35148
rect 16132 35136 16160 35244
rect 16206 35164 16212 35216
rect 16264 35164 16270 35216
rect 12952 35108 16160 35136
rect 12952 35096 12958 35108
rect 6822 35028 6828 35080
rect 6880 35068 6886 35080
rect 13998 35068 14004 35080
rect 6880 35040 14004 35068
rect 6880 35028 6886 35040
rect 13998 35028 14004 35040
rect 14056 35028 14062 35080
rect 14737 35071 14795 35077
rect 14737 35037 14749 35071
rect 14783 35068 14795 35071
rect 14826 35068 14832 35080
rect 14783 35040 14832 35068
rect 14783 35037 14795 35040
rect 14737 35031 14795 35037
rect 14826 35028 14832 35040
rect 14884 35028 14890 35080
rect 15396 35077 15424 35108
rect 15381 35071 15439 35077
rect 15381 35037 15393 35071
rect 15427 35037 15439 35071
rect 15381 35031 15439 35037
rect 15565 35071 15623 35077
rect 15565 35037 15577 35071
rect 15611 35068 15623 35071
rect 15654 35068 15660 35080
rect 15611 35040 15660 35068
rect 15611 35037 15623 35040
rect 15565 35031 15623 35037
rect 15654 35028 15660 35040
rect 15712 35068 15718 35080
rect 16224 35077 16252 35164
rect 16408 35148 16436 35244
rect 19334 35232 19340 35244
rect 19392 35232 19398 35284
rect 23658 35232 23664 35284
rect 23716 35272 23722 35284
rect 25314 35272 25320 35284
rect 23716 35244 25320 35272
rect 23716 35232 23722 35244
rect 25314 35232 25320 35244
rect 25372 35232 25378 35284
rect 26142 35232 26148 35284
rect 26200 35272 26206 35284
rect 26697 35275 26755 35281
rect 26697 35272 26709 35275
rect 26200 35244 26709 35272
rect 26200 35232 26206 35244
rect 26697 35241 26709 35244
rect 26743 35241 26755 35275
rect 27890 35272 27896 35284
rect 27851 35244 27896 35272
rect 26697 35235 26755 35241
rect 27890 35232 27896 35244
rect 27948 35232 27954 35284
rect 16482 35164 16488 35216
rect 16540 35204 16546 35216
rect 16540 35164 16574 35204
rect 16666 35164 16672 35216
rect 16724 35204 16730 35216
rect 20622 35204 20628 35216
rect 16724 35176 20628 35204
rect 16724 35164 16730 35176
rect 20622 35164 20628 35176
rect 20680 35164 20686 35216
rect 22738 35204 22744 35216
rect 22651 35176 22744 35204
rect 22738 35164 22744 35176
rect 22796 35204 22802 35216
rect 23014 35204 23020 35216
rect 22796 35176 23020 35204
rect 22796 35164 22802 35176
rect 23014 35164 23020 35176
rect 23072 35204 23078 35216
rect 25222 35204 25228 35216
rect 23072 35176 25228 35204
rect 23072 35164 23078 35176
rect 25222 35164 25228 35176
rect 25280 35164 25286 35216
rect 25406 35164 25412 35216
rect 25464 35204 25470 35216
rect 25869 35207 25927 35213
rect 25869 35204 25881 35207
rect 25464 35176 25881 35204
rect 25464 35164 25470 35176
rect 25869 35173 25881 35176
rect 25915 35204 25927 35207
rect 27706 35204 27712 35216
rect 25915 35176 27712 35204
rect 25915 35173 25927 35176
rect 25869 35167 25927 35173
rect 27706 35164 27712 35176
rect 27764 35164 27770 35216
rect 31386 35204 31392 35216
rect 31347 35176 31392 35204
rect 31386 35164 31392 35176
rect 31444 35164 31450 35216
rect 16390 35136 16396 35148
rect 16303 35108 16396 35136
rect 16390 35096 16396 35108
rect 16448 35096 16454 35148
rect 16546 35136 16574 35164
rect 17221 35139 17279 35145
rect 16546 35108 16620 35136
rect 16209 35071 16267 35077
rect 15712 35040 16160 35068
rect 15712 35028 15718 35040
rect 10134 34960 10140 35012
rect 10192 35000 10198 35012
rect 12434 35000 12440 35012
rect 10192 34972 12440 35000
rect 10192 34960 10198 34972
rect 12434 34960 12440 34972
rect 12492 34960 12498 35012
rect 14461 35003 14519 35009
rect 14461 34969 14473 35003
rect 14507 35000 14519 35003
rect 16132 35000 16160 35040
rect 16209 35037 16221 35071
rect 16255 35037 16267 35071
rect 16209 35031 16267 35037
rect 16301 35071 16359 35077
rect 16301 35037 16313 35071
rect 16347 35037 16359 35071
rect 16301 35031 16359 35037
rect 16485 35071 16543 35077
rect 16485 35037 16497 35071
rect 16531 35068 16543 35071
rect 16592 35068 16620 35108
rect 17221 35105 17233 35139
rect 17267 35136 17279 35139
rect 29086 35136 29092 35148
rect 17267 35108 29092 35136
rect 17267 35105 17279 35108
rect 17221 35099 17279 35105
rect 16531 35040 16620 35068
rect 16669 35071 16727 35077
rect 16531 35037 16543 35040
rect 16485 35031 16543 35037
rect 16669 35037 16681 35071
rect 16715 35068 16727 35071
rect 16758 35068 16764 35080
rect 16715 35040 16764 35068
rect 16715 35037 16727 35040
rect 16669 35031 16727 35037
rect 16316 35000 16344 35031
rect 16758 35028 16764 35040
rect 16816 35028 16822 35080
rect 17236 35000 17264 35099
rect 29086 35096 29092 35108
rect 29144 35096 29150 35148
rect 19794 35068 19800 35080
rect 19755 35040 19800 35068
rect 19794 35028 19800 35040
rect 19852 35028 19858 35080
rect 20622 35028 20628 35080
rect 20680 35068 20686 35080
rect 20993 35071 21051 35077
rect 20993 35068 21005 35071
rect 20680 35040 21005 35068
rect 20680 35028 20686 35040
rect 20993 35037 21005 35040
rect 21039 35037 21051 35071
rect 20993 35031 21051 35037
rect 21266 35028 21272 35080
rect 21324 35068 21330 35080
rect 23201 35071 23259 35077
rect 23201 35068 23213 35071
rect 21324 35040 23213 35068
rect 21324 35028 21330 35040
rect 23201 35037 23213 35040
rect 23247 35037 23259 35071
rect 23201 35031 23259 35037
rect 23845 35071 23903 35077
rect 23845 35037 23857 35071
rect 23891 35068 23903 35071
rect 24486 35068 24492 35080
rect 23891 35040 24492 35068
rect 23891 35037 23903 35040
rect 23845 35031 23903 35037
rect 24486 35028 24492 35040
rect 24544 35068 24550 35080
rect 24673 35071 24731 35077
rect 24673 35068 24685 35071
rect 24544 35040 24685 35068
rect 24544 35028 24550 35040
rect 24673 35037 24685 35040
rect 24719 35037 24731 35071
rect 24673 35031 24731 35037
rect 24946 35028 24952 35080
rect 25004 35068 25010 35080
rect 25317 35071 25375 35077
rect 25317 35068 25329 35071
rect 25004 35040 25329 35068
rect 25004 35028 25010 35040
rect 25317 35037 25329 35040
rect 25363 35037 25375 35071
rect 25317 35031 25375 35037
rect 26602 35028 26608 35080
rect 26660 35068 26666 35080
rect 26881 35071 26939 35077
rect 26881 35068 26893 35071
rect 26660 35040 26893 35068
rect 26660 35028 26666 35040
rect 26881 35037 26893 35040
rect 26927 35068 26939 35071
rect 27341 35071 27399 35077
rect 27341 35068 27353 35071
rect 26927 35040 27353 35068
rect 26927 35037 26939 35040
rect 26881 35031 26939 35037
rect 27341 35037 27353 35040
rect 27387 35037 27399 35071
rect 30006 35068 30012 35080
rect 29967 35040 30012 35068
rect 27341 35031 27399 35037
rect 30006 35028 30012 35040
rect 30064 35028 30070 35080
rect 33502 35068 33508 35080
rect 33463 35040 33508 35068
rect 33502 35028 33508 35040
rect 33560 35068 33566 35080
rect 33778 35068 33784 35080
rect 33560 35040 33784 35068
rect 33560 35028 33566 35040
rect 33778 35028 33784 35040
rect 33836 35028 33842 35080
rect 34054 35068 34060 35080
rect 33967 35040 34060 35068
rect 34054 35028 34060 35040
rect 34112 35068 34118 35080
rect 36078 35068 36084 35080
rect 34112 35040 35940 35068
rect 36039 35040 36084 35068
rect 34112 35028 34118 35040
rect 14507 34972 16068 35000
rect 16132 34972 17264 35000
rect 14507 34969 14519 34972
rect 14461 34963 14519 34969
rect 14752 34944 14780 34972
rect 9674 34892 9680 34944
rect 9732 34932 9738 34944
rect 11698 34932 11704 34944
rect 9732 34904 11704 34932
rect 9732 34892 9738 34904
rect 11698 34892 11704 34904
rect 11756 34932 11762 34944
rect 12158 34932 12164 34944
rect 11756 34904 12164 34932
rect 11756 34892 11762 34904
rect 12158 34892 12164 34904
rect 12216 34932 12222 34944
rect 12345 34935 12403 34941
rect 12345 34932 12357 34935
rect 12216 34904 12357 34932
rect 12216 34892 12222 34904
rect 12345 34901 12357 34904
rect 12391 34901 12403 34935
rect 14642 34932 14648 34944
rect 14603 34904 14648 34932
rect 12345 34895 12403 34901
rect 14642 34892 14648 34904
rect 14700 34892 14706 34944
rect 14734 34892 14740 34944
rect 14792 34892 14798 34944
rect 16040 34941 16068 34972
rect 22002 34960 22008 35012
rect 22060 35000 22066 35012
rect 30254 35003 30312 35009
rect 30254 35000 30266 35003
rect 22060 34972 30266 35000
rect 22060 34960 22066 34972
rect 30254 34969 30266 34972
rect 30300 34969 30312 35003
rect 30254 34963 30312 34969
rect 31938 34960 31944 35012
rect 31996 35000 32002 35012
rect 33238 35003 33296 35009
rect 33238 35000 33250 35003
rect 31996 34972 33250 35000
rect 31996 34960 32002 34972
rect 33238 34969 33250 34972
rect 33284 34969 33296 35003
rect 33238 34963 33296 34969
rect 34514 34960 34520 35012
rect 34572 35000 34578 35012
rect 35814 35003 35872 35009
rect 35814 35000 35826 35003
rect 34572 34972 35826 35000
rect 34572 34960 34578 34972
rect 35814 34969 35826 34972
rect 35860 34969 35872 35003
rect 35814 34963 35872 34969
rect 16025 34935 16083 34941
rect 16025 34901 16037 34935
rect 16071 34901 16083 34935
rect 19978 34932 19984 34944
rect 19939 34904 19984 34932
rect 16025 34895 16083 34901
rect 19978 34892 19984 34904
rect 20036 34892 20042 34944
rect 20714 34892 20720 34944
rect 20772 34932 20778 34944
rect 21085 34935 21143 34941
rect 21085 34932 21097 34935
rect 20772 34904 21097 34932
rect 20772 34892 20778 34904
rect 21085 34901 21097 34904
rect 21131 34901 21143 34935
rect 21085 34895 21143 34901
rect 21634 34892 21640 34944
rect 21692 34932 21698 34944
rect 21821 34935 21879 34941
rect 21821 34932 21833 34935
rect 21692 34904 21833 34932
rect 21692 34892 21698 34904
rect 21821 34901 21833 34904
rect 21867 34901 21879 34935
rect 21821 34895 21879 34901
rect 22278 34892 22284 34944
rect 22336 34932 22342 34944
rect 23382 34932 23388 34944
rect 22336 34904 23388 34932
rect 22336 34892 22342 34904
rect 23382 34892 23388 34904
rect 23440 34892 23446 34944
rect 24486 34932 24492 34944
rect 24447 34904 24492 34932
rect 24486 34892 24492 34904
rect 24544 34892 24550 34944
rect 25130 34932 25136 34944
rect 25091 34904 25136 34932
rect 25130 34892 25136 34904
rect 25188 34892 25194 34944
rect 28166 34892 28172 34944
rect 28224 34932 28230 34944
rect 28445 34935 28503 34941
rect 28445 34932 28457 34935
rect 28224 34904 28457 34932
rect 28224 34892 28230 34904
rect 28445 34901 28457 34904
rect 28491 34901 28503 34935
rect 28445 34895 28503 34901
rect 31294 34892 31300 34944
rect 31352 34932 31358 34944
rect 32125 34935 32183 34941
rect 32125 34932 32137 34935
rect 31352 34904 32137 34932
rect 31352 34892 31358 34904
rect 32125 34901 32137 34904
rect 32171 34901 32183 34935
rect 32125 34895 32183 34901
rect 34606 34892 34612 34944
rect 34664 34932 34670 34944
rect 34701 34935 34759 34941
rect 34701 34932 34713 34935
rect 34664 34904 34713 34932
rect 34664 34892 34670 34904
rect 34701 34901 34713 34904
rect 34747 34901 34759 34935
rect 35912 34932 35940 35040
rect 36078 35028 36084 35040
rect 36136 35068 36142 35080
rect 36725 35071 36783 35077
rect 36725 35068 36737 35071
rect 36136 35040 36737 35068
rect 36136 35028 36142 35040
rect 36725 35037 36737 35040
rect 36771 35037 36783 35071
rect 36725 35031 36783 35037
rect 36992 35003 37050 35009
rect 36992 34969 37004 35003
rect 37038 35000 37050 35003
rect 37826 35000 37832 35012
rect 37038 34972 37832 35000
rect 37038 34969 37050 34972
rect 36992 34963 37050 34969
rect 37826 34960 37832 34972
rect 37884 34960 37890 35012
rect 36722 34932 36728 34944
rect 35912 34904 36728 34932
rect 34701 34895 34759 34901
rect 36722 34892 36728 34904
rect 36780 34892 36786 34944
rect 37642 34892 37648 34944
rect 37700 34932 37706 34944
rect 38105 34935 38163 34941
rect 38105 34932 38117 34935
rect 37700 34904 38117 34932
rect 37700 34892 37706 34904
rect 38105 34901 38117 34904
rect 38151 34901 38163 34935
rect 38105 34895 38163 34901
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 9398 34688 9404 34740
rect 9456 34728 9462 34740
rect 9585 34731 9643 34737
rect 9585 34728 9597 34731
rect 9456 34700 9597 34728
rect 9456 34688 9462 34700
rect 9585 34697 9597 34700
rect 9631 34728 9643 34731
rect 10870 34728 10876 34740
rect 9631 34700 10876 34728
rect 9631 34697 9643 34700
rect 9585 34691 9643 34697
rect 10870 34688 10876 34700
rect 10928 34688 10934 34740
rect 12075 34731 12133 34737
rect 12075 34697 12087 34731
rect 12121 34728 12133 34731
rect 13538 34728 13544 34740
rect 12121 34700 13544 34728
rect 12121 34697 12133 34700
rect 12075 34691 12133 34697
rect 13538 34688 13544 34700
rect 13596 34688 13602 34740
rect 13722 34688 13728 34740
rect 13780 34728 13786 34740
rect 14553 34731 14611 34737
rect 14553 34728 14565 34731
rect 13780 34700 14565 34728
rect 13780 34688 13786 34700
rect 14553 34697 14565 34700
rect 14599 34697 14611 34731
rect 14553 34691 14611 34697
rect 9950 34620 9956 34672
rect 10008 34660 10014 34672
rect 10045 34663 10103 34669
rect 10045 34660 10057 34663
rect 10008 34632 10057 34660
rect 10008 34620 10014 34632
rect 10045 34629 10057 34632
rect 10091 34660 10103 34663
rect 11882 34660 11888 34672
rect 10091 34632 11888 34660
rect 10091 34629 10103 34632
rect 10045 34623 10103 34629
rect 11882 34620 11888 34632
rect 11940 34660 11946 34672
rect 11940 34632 13584 34660
rect 11940 34620 11946 34632
rect 10226 34592 10232 34604
rect 10187 34564 10232 34592
rect 10226 34552 10232 34564
rect 10284 34552 10290 34604
rect 10318 34552 10324 34604
rect 10376 34592 10382 34604
rect 11977 34595 12035 34601
rect 10376 34564 10421 34592
rect 10376 34552 10382 34564
rect 11977 34561 11989 34595
rect 12023 34561 12035 34595
rect 12158 34592 12164 34604
rect 12119 34564 12164 34592
rect 11977 34555 12035 34561
rect 10134 34524 10140 34536
rect 10060 34496 10140 34524
rect 10060 34465 10088 34496
rect 10134 34484 10140 34496
rect 10192 34484 10198 34536
rect 11992 34524 12020 34555
rect 12158 34552 12164 34564
rect 12216 34552 12222 34604
rect 12253 34595 12311 34601
rect 12253 34561 12265 34595
rect 12299 34592 12311 34595
rect 12342 34592 12348 34604
rect 12299 34564 12348 34592
rect 12299 34561 12311 34564
rect 12253 34555 12311 34561
rect 12342 34552 12348 34564
rect 12400 34552 12406 34604
rect 12894 34592 12900 34604
rect 12855 34564 12900 34592
rect 12894 34552 12900 34564
rect 12952 34552 12958 34604
rect 13556 34601 13584 34632
rect 13081 34595 13139 34601
rect 13081 34561 13093 34595
rect 13127 34561 13139 34595
rect 13081 34555 13139 34561
rect 13541 34595 13599 34601
rect 13541 34561 13553 34595
rect 13587 34561 13599 34595
rect 13541 34555 13599 34561
rect 12802 34524 12808 34536
rect 11992 34496 12808 34524
rect 12802 34484 12808 34496
rect 12860 34484 12866 34536
rect 13096 34468 13124 34555
rect 13633 34527 13691 34533
rect 13633 34493 13645 34527
rect 13679 34524 13691 34527
rect 14090 34524 14096 34536
rect 13679 34496 14096 34524
rect 13679 34493 13691 34496
rect 13633 34487 13691 34493
rect 14090 34484 14096 34496
rect 14148 34484 14154 34536
rect 14568 34524 14596 34691
rect 14642 34688 14648 34740
rect 14700 34728 14706 34740
rect 15010 34728 15016 34740
rect 14700 34700 15016 34728
rect 14700 34688 14706 34700
rect 15010 34688 15016 34700
rect 15068 34728 15074 34740
rect 20993 34731 21051 34737
rect 15068 34700 16574 34728
rect 15068 34688 15074 34700
rect 14734 34660 14740 34672
rect 14695 34632 14740 34660
rect 14734 34620 14740 34632
rect 14792 34620 14798 34672
rect 15654 34660 15660 34672
rect 15615 34632 15660 34660
rect 15654 34620 15660 34632
rect 15712 34620 15718 34672
rect 16546 34660 16574 34700
rect 20993 34697 21005 34731
rect 21039 34697 21051 34731
rect 22002 34728 22008 34740
rect 21963 34700 22008 34728
rect 20993 34691 21051 34697
rect 20438 34660 20444 34672
rect 16546 34632 20444 34660
rect 20438 34620 20444 34632
rect 20496 34620 20502 34672
rect 20714 34660 20720 34672
rect 20548 34632 20720 34660
rect 14918 34592 14924 34604
rect 14879 34564 14924 34592
rect 14918 34552 14924 34564
rect 14976 34552 14982 34604
rect 20548 34592 20576 34632
rect 20714 34620 20720 34632
rect 20772 34620 20778 34672
rect 20456 34564 20576 34592
rect 20625 34595 20683 34601
rect 15194 34524 15200 34536
rect 14568 34496 15200 34524
rect 15194 34484 15200 34496
rect 15252 34484 15258 34536
rect 19426 34484 19432 34536
rect 19484 34524 19490 34536
rect 19613 34527 19671 34533
rect 19613 34524 19625 34527
rect 19484 34496 19625 34524
rect 19484 34484 19490 34496
rect 19613 34493 19625 34496
rect 19659 34524 19671 34527
rect 20254 34524 20260 34536
rect 19659 34496 20260 34524
rect 19659 34493 19671 34496
rect 19613 34487 19671 34493
rect 20254 34484 20260 34496
rect 20312 34484 20318 34536
rect 20456 34533 20484 34564
rect 20625 34561 20637 34595
rect 20671 34561 20683 34595
rect 21008 34592 21036 34691
rect 22002 34688 22008 34700
rect 22060 34688 22066 34740
rect 22741 34731 22799 34737
rect 22741 34697 22753 34731
rect 22787 34697 22799 34731
rect 23382 34728 23388 34740
rect 23343 34700 23388 34728
rect 22741 34691 22799 34697
rect 22756 34660 22784 34691
rect 23382 34688 23388 34700
rect 23440 34688 23446 34740
rect 24302 34728 24308 34740
rect 24263 34700 24308 34728
rect 24302 34688 24308 34700
rect 24360 34688 24366 34740
rect 26234 34728 26240 34740
rect 26195 34700 26240 34728
rect 26234 34688 26240 34700
rect 26292 34688 26298 34740
rect 26970 34728 26976 34740
rect 26931 34700 26976 34728
rect 26970 34688 26976 34700
rect 27028 34688 27034 34740
rect 29086 34728 29092 34740
rect 29047 34700 29092 34728
rect 29086 34688 29092 34700
rect 29144 34688 29150 34740
rect 29178 34688 29184 34740
rect 29236 34728 29242 34740
rect 29236 34700 31754 34728
rect 29236 34688 29242 34700
rect 27982 34660 27988 34672
rect 22756 34632 27988 34660
rect 27982 34620 27988 34632
rect 28040 34620 28046 34672
rect 29638 34620 29644 34672
rect 29696 34660 29702 34672
rect 30006 34660 30012 34672
rect 29696 34632 30012 34660
rect 29696 34620 29702 34632
rect 30006 34620 30012 34632
rect 30064 34660 30070 34672
rect 31726 34660 31754 34700
rect 34158 34663 34216 34669
rect 34158 34660 34170 34663
rect 30064 34632 30512 34660
rect 31726 34632 34170 34660
rect 30064 34620 30070 34632
rect 21821 34595 21879 34601
rect 21821 34592 21833 34595
rect 21008 34564 21833 34592
rect 20625 34555 20683 34561
rect 21821 34561 21833 34564
rect 21867 34561 21879 34595
rect 22554 34592 22560 34604
rect 22515 34564 22560 34592
rect 21821 34555 21879 34561
rect 20441 34527 20499 34533
rect 20441 34493 20453 34527
rect 20487 34493 20499 34527
rect 20441 34487 20499 34493
rect 20533 34527 20591 34533
rect 20533 34493 20545 34527
rect 20579 34493 20591 34527
rect 20640 34524 20668 34555
rect 22554 34552 22560 34564
rect 22612 34552 22618 34604
rect 23198 34592 23204 34604
rect 23159 34564 23204 34592
rect 23198 34552 23204 34564
rect 23256 34552 23262 34604
rect 24854 34552 24860 34604
rect 24912 34592 24918 34604
rect 25418 34595 25476 34601
rect 25418 34592 25430 34595
rect 24912 34564 25430 34592
rect 24912 34552 24918 34564
rect 25418 34561 25430 34564
rect 25464 34561 25476 34595
rect 25418 34555 25476 34561
rect 25590 34552 25596 34604
rect 25648 34592 25654 34604
rect 25685 34595 25743 34601
rect 25685 34592 25697 34595
rect 25648 34564 25697 34592
rect 25648 34552 25654 34564
rect 25685 34561 25697 34564
rect 25731 34561 25743 34595
rect 28074 34592 28080 34604
rect 28132 34601 28138 34604
rect 28044 34564 28080 34592
rect 25685 34555 25743 34561
rect 28074 34552 28080 34564
rect 28132 34555 28144 34601
rect 28353 34595 28411 34601
rect 28353 34561 28365 34595
rect 28399 34592 28411 34595
rect 29656 34592 29684 34620
rect 28399 34564 29684 34592
rect 28399 34561 28411 34564
rect 28353 34555 28411 34561
rect 28132 34552 28138 34555
rect 30190 34552 30196 34604
rect 30248 34601 30254 34604
rect 30484 34601 30512 34632
rect 34158 34629 34170 34632
rect 34204 34629 34216 34663
rect 34158 34623 34216 34629
rect 30248 34592 30260 34601
rect 30469 34595 30527 34601
rect 30248 34564 30293 34592
rect 30248 34555 30260 34564
rect 30469 34561 30481 34595
rect 30515 34561 30527 34595
rect 30469 34555 30527 34561
rect 30248 34552 30254 34555
rect 34790 34552 34796 34604
rect 34848 34592 34854 34604
rect 38194 34592 38200 34604
rect 34848 34564 38200 34592
rect 34848 34552 34854 34564
rect 38194 34552 38200 34564
rect 38252 34552 38258 34604
rect 21634 34524 21640 34536
rect 20640 34496 21640 34524
rect 20533 34487 20591 34493
rect 10045 34459 10103 34465
rect 10045 34425 10057 34459
rect 10091 34425 10103 34459
rect 13078 34456 13084 34468
rect 12991 34428 13084 34456
rect 10045 34419 10103 34425
rect 13078 34416 13084 34428
rect 13136 34456 13142 34468
rect 14918 34456 14924 34468
rect 13136 34428 14924 34456
rect 13136 34416 13142 34428
rect 14918 34416 14924 34428
rect 14976 34416 14982 34468
rect 20548 34456 20576 34487
rect 21634 34484 21640 34496
rect 21692 34484 21698 34536
rect 34425 34527 34483 34533
rect 34425 34493 34437 34527
rect 34471 34493 34483 34527
rect 34425 34487 34483 34493
rect 35897 34527 35955 34533
rect 35897 34493 35909 34527
rect 35943 34524 35955 34527
rect 35986 34524 35992 34536
rect 35943 34496 35992 34524
rect 35943 34493 35955 34496
rect 35897 34487 35955 34493
rect 20898 34456 20904 34468
rect 20548 34428 20904 34456
rect 20898 34416 20904 34428
rect 20956 34416 20962 34468
rect 12986 34388 12992 34400
rect 12947 34360 12992 34388
rect 12986 34348 12992 34360
rect 13044 34348 13050 34400
rect 16574 34348 16580 34400
rect 16632 34388 16638 34400
rect 16850 34388 16856 34400
rect 16632 34360 16856 34388
rect 16632 34348 16638 34360
rect 16850 34348 16856 34360
rect 16908 34348 16914 34400
rect 33042 34388 33048 34400
rect 33003 34360 33048 34388
rect 33042 34348 33048 34360
rect 33100 34348 33106 34400
rect 33134 34348 33140 34400
rect 33192 34388 33198 34400
rect 33502 34388 33508 34400
rect 33192 34360 33508 34388
rect 33192 34348 33198 34360
rect 33502 34348 33508 34360
rect 33560 34388 33566 34400
rect 34440 34388 34468 34487
rect 35986 34484 35992 34496
rect 36044 34524 36050 34536
rect 37277 34527 37335 34533
rect 37277 34524 37289 34527
rect 36044 34496 37289 34524
rect 36044 34484 36050 34496
rect 37277 34493 37289 34496
rect 37323 34493 37335 34527
rect 37277 34487 37335 34493
rect 36262 34456 36268 34468
rect 36175 34428 36268 34456
rect 36262 34416 36268 34428
rect 36320 34456 36326 34468
rect 37829 34459 37887 34465
rect 37829 34456 37841 34459
rect 36320 34428 37841 34456
rect 36320 34416 36326 34428
rect 37829 34425 37841 34428
rect 37875 34425 37887 34459
rect 37829 34419 37887 34425
rect 36354 34388 36360 34400
rect 33560 34360 34468 34388
rect 36315 34360 36360 34388
rect 33560 34348 33566 34360
rect 36354 34348 36360 34360
rect 36412 34348 36418 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 10318 34144 10324 34196
rect 10376 34184 10382 34196
rect 10597 34187 10655 34193
rect 10597 34184 10609 34187
rect 10376 34156 10609 34184
rect 10376 34144 10382 34156
rect 10597 34153 10609 34156
rect 10643 34153 10655 34187
rect 10597 34147 10655 34153
rect 11716 34156 12434 34184
rect 11716 34057 11744 34156
rect 12250 34116 12256 34128
rect 12211 34088 12256 34116
rect 12250 34076 12256 34088
rect 12308 34076 12314 34128
rect 12406 34116 12434 34156
rect 15102 34144 15108 34196
rect 15160 34184 15166 34196
rect 15197 34187 15255 34193
rect 15197 34184 15209 34187
rect 15160 34156 15209 34184
rect 15160 34144 15166 34156
rect 15197 34153 15209 34156
rect 15243 34153 15255 34187
rect 15197 34147 15255 34153
rect 16666 34144 16672 34196
rect 16724 34184 16730 34196
rect 22186 34184 22192 34196
rect 16724 34156 16769 34184
rect 22147 34156 22192 34184
rect 16724 34144 16730 34156
rect 22186 34144 22192 34156
rect 22244 34144 22250 34196
rect 22925 34187 22983 34193
rect 22925 34153 22937 34187
rect 22971 34184 22983 34187
rect 23198 34184 23204 34196
rect 22971 34156 23204 34184
rect 22971 34153 22983 34156
rect 22925 34147 22983 34153
rect 23198 34144 23204 34156
rect 23256 34144 23262 34196
rect 24946 34184 24952 34196
rect 24907 34156 24952 34184
rect 24946 34144 24952 34156
rect 25004 34144 25010 34196
rect 25406 34144 25412 34196
rect 25464 34184 25470 34196
rect 25593 34187 25651 34193
rect 25593 34184 25605 34187
rect 25464 34156 25605 34184
rect 25464 34144 25470 34156
rect 25593 34153 25605 34156
rect 25639 34184 25651 34187
rect 25774 34184 25780 34196
rect 25639 34156 25780 34184
rect 25639 34153 25651 34156
rect 25593 34147 25651 34153
rect 25774 34144 25780 34156
rect 25832 34144 25838 34196
rect 28994 34184 29000 34196
rect 28955 34156 29000 34184
rect 28994 34144 29000 34156
rect 29052 34184 29058 34196
rect 30190 34184 30196 34196
rect 29052 34156 30196 34184
rect 29052 34144 29058 34156
rect 30190 34144 30196 34156
rect 30248 34144 30254 34196
rect 35986 34184 35992 34196
rect 31726 34156 35992 34184
rect 12805 34119 12863 34125
rect 12805 34116 12817 34119
rect 12406 34088 12817 34116
rect 12805 34085 12817 34088
rect 12851 34085 12863 34119
rect 12805 34079 12863 34085
rect 16390 34076 16396 34128
rect 16448 34116 16454 34128
rect 26697 34119 26755 34125
rect 26697 34116 26709 34119
rect 16448 34088 26709 34116
rect 16448 34076 16454 34088
rect 26697 34085 26709 34088
rect 26743 34085 26755 34119
rect 26697 34079 26755 34085
rect 10045 34051 10103 34057
rect 10045 34017 10057 34051
rect 10091 34048 10103 34051
rect 11701 34051 11759 34057
rect 11701 34048 11713 34051
rect 10091 34020 11713 34048
rect 10091 34017 10103 34020
rect 10045 34011 10103 34017
rect 11701 34017 11713 34020
rect 11747 34017 11759 34051
rect 11701 34011 11759 34017
rect 11977 34051 12035 34057
rect 11977 34017 11989 34051
rect 12023 34048 12035 34051
rect 12986 34048 12992 34060
rect 12023 34020 12992 34048
rect 12023 34017 12035 34020
rect 11977 34011 12035 34017
rect 12986 34008 12992 34020
rect 13044 34008 13050 34060
rect 14918 34008 14924 34060
rect 14976 34048 14982 34060
rect 20901 34051 20959 34057
rect 14976 34020 17816 34048
rect 14976 34008 14982 34020
rect 9214 33980 9220 33992
rect 9175 33952 9220 33980
rect 9214 33940 9220 33952
rect 9272 33940 9278 33992
rect 9398 33980 9404 33992
rect 9359 33952 9404 33980
rect 9398 33940 9404 33952
rect 9456 33980 9462 33992
rect 9456 33952 10180 33980
rect 9456 33940 9462 33952
rect 10152 33912 10180 33952
rect 10226 33940 10232 33992
rect 10284 33980 10290 33992
rect 11517 33983 11575 33989
rect 11517 33980 11529 33983
rect 10284 33952 11529 33980
rect 10284 33940 10290 33952
rect 11517 33949 11529 33952
rect 11563 33949 11575 33983
rect 11517 33943 11575 33949
rect 11882 33940 11888 33992
rect 11940 33980 11946 33992
rect 12253 33983 12311 33989
rect 12253 33980 12265 33983
rect 11940 33952 12265 33980
rect 11940 33940 11946 33952
rect 12253 33949 12265 33952
rect 12299 33949 12311 33983
rect 12253 33943 12311 33949
rect 13173 33983 13231 33989
rect 13173 33949 13185 33983
rect 13219 33980 13231 33983
rect 13814 33980 13820 33992
rect 13219 33952 13820 33980
rect 13219 33949 13231 33952
rect 13173 33943 13231 33949
rect 13814 33940 13820 33952
rect 13872 33940 13878 33992
rect 14090 33980 14096 33992
rect 14051 33952 14096 33980
rect 14090 33940 14096 33952
rect 14148 33940 14154 33992
rect 17678 33980 17684 33992
rect 14292 33952 17684 33980
rect 10152 33884 10364 33912
rect 9401 33847 9459 33853
rect 9401 33813 9413 33847
rect 9447 33844 9459 33847
rect 10137 33847 10195 33853
rect 10137 33844 10149 33847
rect 9447 33816 10149 33844
rect 9447 33813 9459 33816
rect 9401 33807 9459 33813
rect 10137 33813 10149 33816
rect 10183 33813 10195 33847
rect 10137 33807 10195 33813
rect 10229 33847 10287 33853
rect 10229 33813 10241 33847
rect 10275 33844 10287 33847
rect 10336 33844 10364 33884
rect 12894 33872 12900 33924
rect 12952 33912 12958 33924
rect 12989 33915 13047 33921
rect 12989 33912 13001 33915
rect 12952 33884 13001 33912
rect 12952 33872 12958 33884
rect 12989 33881 13001 33884
rect 13035 33881 13047 33915
rect 12989 33875 13047 33881
rect 14292 33853 14320 33952
rect 17678 33940 17684 33952
rect 17736 33940 17742 33992
rect 17788 33980 17816 34020
rect 20901 34017 20913 34051
rect 20947 34048 20959 34051
rect 22094 34048 22100 34060
rect 20947 34020 22100 34048
rect 20947 34017 20959 34020
rect 20901 34011 20959 34017
rect 22094 34008 22100 34020
rect 22152 34008 22158 34060
rect 23198 34008 23204 34060
rect 23256 34048 23262 34060
rect 23477 34051 23535 34057
rect 23477 34048 23489 34051
rect 23256 34020 23489 34048
rect 23256 34008 23262 34020
rect 23477 34017 23489 34020
rect 23523 34017 23535 34051
rect 23477 34011 23535 34017
rect 24489 34051 24547 34057
rect 24489 34017 24501 34051
rect 24535 34048 24547 34051
rect 24578 34048 24584 34060
rect 24535 34020 24584 34048
rect 24535 34017 24547 34020
rect 24489 34011 24547 34017
rect 24578 34008 24584 34020
rect 24636 34008 24642 34060
rect 24762 34008 24768 34060
rect 24820 34048 24826 34060
rect 26053 34051 26111 34057
rect 26053 34048 26065 34051
rect 24820 34020 26065 34048
rect 24820 34008 24826 34020
rect 26053 34017 26065 34020
rect 26099 34017 26111 34051
rect 26053 34011 26111 34017
rect 28077 34051 28135 34057
rect 28077 34017 28089 34051
rect 28123 34048 28135 34051
rect 29638 34048 29644 34060
rect 28123 34020 29644 34048
rect 28123 34017 28135 34020
rect 28077 34011 28135 34017
rect 29638 34008 29644 34020
rect 29696 34008 29702 34060
rect 17844 33983 17902 33989
rect 18049 33983 18107 33989
rect 17844 33980 17856 33983
rect 17788 33952 17856 33980
rect 17844 33949 17856 33952
rect 17890 33949 17902 33983
rect 17844 33943 17902 33949
rect 17944 33977 18002 33983
rect 17944 33943 17956 33977
rect 17990 33943 18002 33977
rect 18049 33949 18061 33983
rect 18095 33980 18107 33983
rect 18095 33952 19380 33980
rect 18095 33949 18107 33952
rect 18049 33943 18107 33949
rect 17944 33937 18002 33943
rect 15010 33912 15016 33924
rect 14971 33884 15016 33912
rect 15010 33872 15016 33884
rect 15068 33872 15074 33924
rect 15194 33872 15200 33924
rect 15252 33921 15258 33924
rect 15252 33915 15271 33921
rect 15259 33881 15271 33915
rect 15252 33875 15271 33881
rect 16393 33915 16451 33921
rect 16393 33881 16405 33915
rect 16439 33912 16451 33915
rect 16482 33912 16488 33924
rect 16439 33884 16488 33912
rect 16439 33881 16451 33884
rect 16393 33875 16451 33881
rect 15252 33872 15258 33875
rect 16482 33872 16488 33884
rect 16540 33872 16546 33924
rect 16574 33872 16580 33924
rect 16632 33912 16638 33924
rect 16632 33884 16677 33912
rect 16632 33872 16638 33884
rect 10275 33816 10364 33844
rect 14277 33847 14335 33853
rect 10275 33813 10287 33816
rect 10229 33807 10287 33813
rect 14277 33813 14289 33847
rect 14323 33813 14335 33847
rect 14277 33807 14335 33813
rect 15381 33847 15439 33853
rect 15381 33813 15393 33847
rect 15427 33844 15439 33847
rect 16666 33844 16672 33856
rect 15427 33816 16672 33844
rect 15427 33813 15439 33816
rect 15381 33807 15439 33813
rect 16666 33804 16672 33816
rect 16724 33804 16730 33856
rect 17972 33844 18000 33937
rect 18322 33912 18328 33924
rect 18283 33884 18328 33912
rect 18322 33872 18328 33884
rect 18380 33872 18386 33924
rect 19352 33921 19380 33952
rect 20438 33940 20444 33992
rect 20496 33980 20502 33992
rect 21361 33983 21419 33989
rect 21361 33980 21373 33983
rect 20496 33952 21373 33980
rect 20496 33940 20502 33952
rect 21361 33949 21373 33952
rect 21407 33949 21419 33983
rect 21361 33943 21419 33949
rect 21818 33940 21824 33992
rect 21876 33980 21882 33992
rect 22005 33983 22063 33989
rect 22005 33980 22017 33983
rect 21876 33952 22017 33980
rect 21876 33940 21882 33952
rect 22005 33949 22017 33952
rect 22051 33949 22063 33983
rect 22005 33943 22063 33949
rect 23385 33983 23443 33989
rect 23385 33949 23397 33983
rect 23431 33980 23443 33983
rect 25130 33980 25136 33992
rect 23431 33952 25136 33980
rect 23431 33949 23443 33952
rect 23385 33943 23443 33949
rect 25130 33940 25136 33952
rect 25188 33940 25194 33992
rect 27798 33980 27804 33992
rect 27856 33989 27862 33992
rect 27768 33952 27804 33980
rect 27798 33940 27804 33952
rect 27856 33943 27868 33989
rect 27856 33940 27862 33943
rect 19337 33915 19395 33921
rect 19337 33881 19349 33915
rect 19383 33912 19395 33915
rect 31726 33912 31754 34156
rect 35986 34144 35992 34156
rect 36044 34184 36050 34196
rect 36081 34187 36139 34193
rect 36081 34184 36093 34187
rect 36044 34156 36093 34184
rect 36044 34144 36050 34156
rect 36081 34153 36093 34156
rect 36127 34153 36139 34187
rect 36081 34147 36139 34153
rect 34701 33983 34759 33989
rect 34701 33949 34713 33983
rect 34747 33980 34759 33983
rect 35894 33980 35900 33992
rect 34747 33952 35900 33980
rect 34747 33949 34759 33952
rect 34701 33943 34759 33949
rect 35894 33940 35900 33952
rect 35952 33980 35958 33992
rect 36078 33980 36084 33992
rect 35952 33952 36084 33980
rect 35952 33940 35958 33952
rect 36078 33940 36084 33952
rect 36136 33980 36142 33992
rect 36725 33983 36783 33989
rect 36725 33980 36737 33983
rect 36136 33952 36737 33980
rect 36136 33940 36142 33952
rect 36725 33949 36737 33952
rect 36771 33949 36783 33983
rect 36725 33943 36783 33949
rect 19383 33884 31754 33912
rect 32953 33915 33011 33921
rect 19383 33881 19395 33884
rect 19337 33875 19395 33881
rect 32953 33881 32965 33915
rect 32999 33912 33011 33915
rect 33226 33912 33232 33924
rect 32999 33884 33232 33912
rect 32999 33881 33011 33884
rect 32953 33875 33011 33881
rect 33226 33872 33232 33884
rect 33284 33872 33290 33924
rect 34514 33872 34520 33924
rect 34572 33912 34578 33924
rect 34946 33915 35004 33921
rect 34946 33912 34958 33915
rect 34572 33884 34958 33912
rect 34572 33872 34578 33884
rect 34946 33881 34958 33884
rect 34992 33881 35004 33915
rect 36992 33915 37050 33921
rect 34946 33875 35004 33881
rect 35866 33884 36216 33912
rect 18046 33844 18052 33856
rect 17972 33816 18052 33844
rect 18046 33804 18052 33816
rect 18104 33804 18110 33856
rect 21545 33847 21603 33853
rect 21545 33813 21557 33847
rect 21591 33844 21603 33847
rect 23106 33844 23112 33856
rect 21591 33816 23112 33844
rect 21591 33813 21603 33816
rect 21545 33807 21603 33813
rect 23106 33804 23112 33816
rect 23164 33804 23170 33856
rect 23293 33847 23351 33853
rect 23293 33813 23305 33847
rect 23339 33844 23351 33847
rect 24026 33844 24032 33856
rect 23339 33816 24032 33844
rect 23339 33813 23351 33816
rect 23293 33807 23351 33813
rect 24026 33804 24032 33816
rect 24084 33844 24090 33856
rect 24578 33844 24584 33856
rect 24084 33816 24584 33844
rect 24084 33804 24090 33816
rect 24578 33804 24584 33816
rect 24636 33804 24642 33856
rect 31665 33847 31723 33853
rect 31665 33813 31677 33847
rect 31711 33844 31723 33847
rect 33134 33844 33140 33856
rect 31711 33816 33140 33844
rect 31711 33813 31723 33816
rect 31665 33807 31723 33813
rect 33134 33804 33140 33816
rect 33192 33804 33198 33856
rect 34238 33804 34244 33856
rect 34296 33844 34302 33856
rect 35866 33844 35894 33884
rect 34296 33816 35894 33844
rect 36188 33844 36216 33884
rect 36992 33881 37004 33915
rect 37038 33912 37050 33915
rect 37090 33912 37096 33924
rect 37038 33884 37096 33912
rect 37038 33881 37050 33884
rect 36992 33875 37050 33881
rect 37090 33872 37096 33884
rect 37148 33872 37154 33924
rect 38105 33847 38163 33853
rect 38105 33844 38117 33847
rect 36188 33816 38117 33844
rect 34296 33804 34302 33816
rect 38105 33813 38117 33816
rect 38151 33813 38163 33847
rect 38105 33807 38163 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 8754 33640 8760 33652
rect 8715 33612 8760 33640
rect 8754 33600 8760 33612
rect 8812 33600 8818 33652
rect 10226 33600 10232 33652
rect 10284 33640 10290 33652
rect 10781 33643 10839 33649
rect 10781 33640 10793 33643
rect 10284 33612 10793 33640
rect 10284 33600 10290 33612
rect 10781 33609 10793 33612
rect 10827 33609 10839 33643
rect 10781 33603 10839 33609
rect 12989 33643 13047 33649
rect 12989 33609 13001 33643
rect 13035 33640 13047 33643
rect 13078 33640 13084 33652
rect 13035 33612 13084 33640
rect 13035 33609 13047 33612
rect 12989 33603 13047 33609
rect 13078 33600 13084 33612
rect 13136 33600 13142 33652
rect 13170 33600 13176 33652
rect 13228 33640 13234 33652
rect 13354 33640 13360 33652
rect 13228 33612 13360 33640
rect 13228 33600 13234 33612
rect 13354 33600 13360 33612
rect 13412 33600 13418 33652
rect 19981 33643 20039 33649
rect 19981 33609 19993 33643
rect 20027 33640 20039 33643
rect 20070 33640 20076 33652
rect 20027 33612 20076 33640
rect 20027 33609 20039 33612
rect 19981 33603 20039 33609
rect 20070 33600 20076 33612
rect 20128 33600 20134 33652
rect 20438 33640 20444 33652
rect 20399 33612 20444 33640
rect 20438 33600 20444 33612
rect 20496 33600 20502 33652
rect 21818 33640 21824 33652
rect 21779 33612 21824 33640
rect 21818 33600 21824 33612
rect 21876 33600 21882 33652
rect 22554 33600 22560 33652
rect 22612 33640 22618 33652
rect 23017 33643 23075 33649
rect 23017 33640 23029 33643
rect 22612 33612 23029 33640
rect 22612 33600 22618 33612
rect 23017 33609 23029 33612
rect 23063 33609 23075 33643
rect 23017 33603 23075 33609
rect 23477 33643 23535 33649
rect 23477 33609 23489 33643
rect 23523 33640 23535 33643
rect 24486 33640 24492 33652
rect 23523 33612 24492 33640
rect 23523 33609 23535 33612
rect 23477 33603 23535 33609
rect 24486 33600 24492 33612
rect 24544 33600 24550 33652
rect 36265 33643 36323 33649
rect 36265 33609 36277 33643
rect 36311 33640 36323 33643
rect 37734 33640 37740 33652
rect 36311 33612 37740 33640
rect 36311 33609 36323 33612
rect 36265 33603 36323 33609
rect 37734 33600 37740 33612
rect 37792 33600 37798 33652
rect 8772 33504 8800 33600
rect 9401 33575 9459 33581
rect 9401 33541 9413 33575
rect 9447 33572 9459 33575
rect 13814 33572 13820 33584
rect 9447 33544 10456 33572
rect 9447 33541 9459 33544
rect 9401 33535 9459 33541
rect 8846 33504 8852 33516
rect 8759 33476 8852 33504
rect 8846 33464 8852 33476
rect 8904 33504 8910 33516
rect 9309 33507 9367 33513
rect 9309 33504 9321 33507
rect 8904 33476 9321 33504
rect 8904 33464 8910 33476
rect 9309 33473 9321 33476
rect 9355 33473 9367 33507
rect 9309 33467 9367 33473
rect 9493 33507 9551 33513
rect 9493 33473 9505 33507
rect 9539 33504 9551 33507
rect 9674 33504 9680 33516
rect 9539 33476 9680 33504
rect 9539 33473 9551 33476
rect 9493 33467 9551 33473
rect 9674 33464 9680 33476
rect 9732 33464 9738 33516
rect 10428 33513 10456 33544
rect 10520 33544 12434 33572
rect 10413 33507 10471 33513
rect 10413 33473 10425 33507
rect 10459 33473 10471 33507
rect 10413 33467 10471 33473
rect 9214 33396 9220 33448
rect 9272 33436 9278 33448
rect 10520 33436 10548 33544
rect 10597 33507 10655 33513
rect 10597 33473 10609 33507
rect 10643 33504 10655 33507
rect 11517 33507 11575 33513
rect 11517 33504 11529 33507
rect 10643 33476 11529 33504
rect 10643 33473 10655 33476
rect 10597 33467 10655 33473
rect 11517 33473 11529 33476
rect 11563 33473 11575 33507
rect 11517 33467 11575 33473
rect 9272 33408 10548 33436
rect 9272 33396 9278 33408
rect 10520 33309 10548 33408
rect 10505 33303 10563 33309
rect 10505 33269 10517 33303
rect 10551 33269 10563 33303
rect 11532 33300 11560 33467
rect 12406 33436 12434 33544
rect 12728 33544 13820 33572
rect 12728 33513 12756 33544
rect 13814 33532 13820 33544
rect 13872 33532 13878 33584
rect 22281 33575 22339 33581
rect 22281 33541 22293 33575
rect 22327 33572 22339 33575
rect 26050 33572 26056 33584
rect 22327 33544 26056 33572
rect 22327 33541 22339 33544
rect 22281 33535 22339 33541
rect 26050 33532 26056 33544
rect 26108 33532 26114 33584
rect 12713 33507 12771 33513
rect 12713 33473 12725 33507
rect 12759 33473 12771 33507
rect 12713 33467 12771 33473
rect 12802 33464 12808 33516
rect 12860 33504 12866 33516
rect 13170 33504 13176 33516
rect 12860 33476 13176 33504
rect 12860 33464 12866 33476
rect 13170 33464 13176 33476
rect 13228 33464 13234 33516
rect 13909 33507 13967 33513
rect 13909 33473 13921 33507
rect 13955 33504 13967 33507
rect 14090 33504 14096 33516
rect 13955 33476 14096 33504
rect 13955 33473 13967 33476
rect 13909 33467 13967 33473
rect 14090 33464 14096 33476
rect 14148 33464 14154 33516
rect 16666 33504 16672 33516
rect 16627 33476 16672 33504
rect 16666 33464 16672 33476
rect 16724 33464 16730 33516
rect 18230 33504 18236 33516
rect 18191 33476 18236 33504
rect 18230 33464 18236 33476
rect 18288 33464 18294 33516
rect 20070 33504 20076 33516
rect 20031 33476 20076 33504
rect 20070 33464 20076 33476
rect 20128 33504 20134 33516
rect 20901 33507 20959 33513
rect 20901 33504 20913 33507
rect 20128 33476 20913 33504
rect 20128 33464 20134 33476
rect 20901 33473 20913 33476
rect 20947 33473 20959 33507
rect 20901 33467 20959 33473
rect 22189 33507 22247 33513
rect 22189 33473 22201 33507
rect 22235 33504 22247 33507
rect 22738 33504 22744 33516
rect 22235 33476 22744 33504
rect 22235 33473 22247 33476
rect 22189 33467 22247 33473
rect 22738 33464 22744 33476
rect 22796 33464 22802 33516
rect 22922 33464 22928 33516
rect 22980 33504 22986 33516
rect 23385 33507 23443 33513
rect 23385 33504 23397 33507
rect 22980 33476 23397 33504
rect 22980 33464 22986 33476
rect 23385 33473 23397 33476
rect 23431 33504 23443 33507
rect 24305 33507 24363 33513
rect 24305 33504 24317 33507
rect 23431 33476 24317 33504
rect 23431 33473 23443 33476
rect 23385 33467 23443 33473
rect 24305 33473 24317 33476
rect 24351 33504 24363 33507
rect 27614 33504 27620 33516
rect 24351 33476 27620 33504
rect 24351 33473 24363 33476
rect 24305 33467 24363 33473
rect 27614 33464 27620 33476
rect 27672 33464 27678 33516
rect 27798 33464 27804 33516
rect 27856 33504 27862 33516
rect 28629 33507 28687 33513
rect 28629 33504 28641 33507
rect 27856 33476 28641 33504
rect 27856 33464 27862 33476
rect 28629 33473 28641 33476
rect 28675 33473 28687 33507
rect 28629 33467 28687 33473
rect 33226 33464 33232 33516
rect 33284 33504 33290 33516
rect 33781 33507 33839 33513
rect 33781 33504 33793 33507
rect 33284 33476 33793 33504
rect 33284 33464 33290 33476
rect 33781 33473 33793 33476
rect 33827 33473 33839 33507
rect 33781 33467 33839 33473
rect 36081 33507 36139 33513
rect 36081 33473 36093 33507
rect 36127 33504 36139 33507
rect 36354 33504 36360 33516
rect 36127 33476 36360 33504
rect 36127 33473 36139 33476
rect 36081 33467 36139 33473
rect 36354 33464 36360 33476
rect 36412 33464 36418 33516
rect 12820 33436 12848 33464
rect 12406 33408 12848 33436
rect 18046 33396 18052 33448
rect 18104 33436 18110 33448
rect 19889 33439 19947 33445
rect 19889 33436 19901 33439
rect 18104 33408 19901 33436
rect 18104 33396 18110 33408
rect 19889 33405 19901 33408
rect 19935 33436 19947 33439
rect 20622 33436 20628 33448
rect 19935 33408 20628 33436
rect 19935 33405 19947 33408
rect 19889 33399 19947 33405
rect 20622 33396 20628 33408
rect 20680 33396 20686 33448
rect 22465 33439 22523 33445
rect 22465 33405 22477 33439
rect 22511 33436 22523 33439
rect 23198 33436 23204 33448
rect 22511 33408 23204 33436
rect 22511 33405 22523 33408
rect 22465 33399 22523 33405
rect 23198 33396 23204 33408
rect 23256 33436 23262 33448
rect 23569 33439 23627 33445
rect 23569 33436 23581 33439
rect 23256 33408 23581 33436
rect 23256 33396 23262 33408
rect 23569 33405 23581 33408
rect 23615 33405 23627 33439
rect 23569 33399 23627 33405
rect 35529 33439 35587 33445
rect 35529 33405 35541 33439
rect 35575 33436 35587 33439
rect 35894 33436 35900 33448
rect 35575 33408 35900 33436
rect 35575 33405 35587 33408
rect 35529 33399 35587 33405
rect 35894 33396 35900 33408
rect 35952 33396 35958 33448
rect 16853 33371 16911 33377
rect 16853 33337 16865 33371
rect 16899 33368 16911 33371
rect 23658 33368 23664 33380
rect 16899 33340 23664 33368
rect 16899 33337 16911 33340
rect 16853 33331 16911 33337
rect 23658 33328 23664 33340
rect 23716 33328 23722 33380
rect 12710 33300 12716 33312
rect 11532 33272 12716 33300
rect 10505 33263 10563 33269
rect 12710 33260 12716 33272
rect 12768 33260 12774 33312
rect 14093 33303 14151 33309
rect 14093 33269 14105 33303
rect 14139 33300 14151 33303
rect 14366 33300 14372 33312
rect 14139 33272 14372 33300
rect 14139 33269 14151 33272
rect 14093 33263 14151 33269
rect 14366 33260 14372 33272
rect 14424 33300 14430 33312
rect 14829 33303 14887 33309
rect 14829 33300 14841 33303
rect 14424 33272 14841 33300
rect 14424 33260 14430 33272
rect 14829 33269 14841 33272
rect 14875 33300 14887 33303
rect 15102 33300 15108 33312
rect 14875 33272 15108 33300
rect 14875 33269 14887 33272
rect 14829 33263 14887 33269
rect 15102 33260 15108 33272
rect 15160 33300 15166 33312
rect 16758 33300 16764 33312
rect 15160 33272 16764 33300
rect 15160 33260 15166 33272
rect 16758 33260 16764 33272
rect 16816 33260 16822 33312
rect 17589 33303 17647 33309
rect 17589 33269 17601 33303
rect 17635 33300 17647 33303
rect 17678 33300 17684 33312
rect 17635 33272 17684 33300
rect 17635 33269 17647 33272
rect 17589 33263 17647 33269
rect 17678 33260 17684 33272
rect 17736 33300 17742 33312
rect 18138 33300 18144 33312
rect 17736 33272 18144 33300
rect 17736 33260 17742 33272
rect 18138 33260 18144 33272
rect 18196 33260 18202 33312
rect 18417 33303 18475 33309
rect 18417 33269 18429 33303
rect 18463 33300 18475 33303
rect 20806 33300 20812 33312
rect 18463 33272 20812 33300
rect 18463 33269 18475 33272
rect 18417 33263 18475 33269
rect 20806 33260 20812 33272
rect 20864 33260 20870 33312
rect 29638 33260 29644 33312
rect 29696 33300 29702 33312
rect 29917 33303 29975 33309
rect 29917 33300 29929 33303
rect 29696 33272 29929 33300
rect 29696 33260 29702 33272
rect 29917 33269 29929 33272
rect 29963 33269 29975 33303
rect 29917 33263 29975 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 9674 33056 9680 33108
rect 9732 33096 9738 33108
rect 9769 33099 9827 33105
rect 9769 33096 9781 33099
rect 9732 33068 9781 33096
rect 9732 33056 9738 33068
rect 9769 33065 9781 33068
rect 9815 33065 9827 33099
rect 9769 33059 9827 33065
rect 12342 33056 12348 33108
rect 12400 33096 12406 33108
rect 12713 33099 12771 33105
rect 12713 33096 12725 33099
rect 12400 33068 12725 33096
rect 12400 33056 12406 33068
rect 12713 33065 12725 33068
rect 12759 33065 12771 33099
rect 12713 33059 12771 33065
rect 18230 33056 18236 33108
rect 18288 33096 18294 33108
rect 18417 33099 18475 33105
rect 18417 33096 18429 33099
rect 18288 33068 18429 33096
rect 18288 33056 18294 33068
rect 18417 33065 18429 33068
rect 18463 33065 18475 33099
rect 18417 33059 18475 33065
rect 22094 33056 22100 33108
rect 22152 33096 22158 33108
rect 28261 33099 28319 33105
rect 28261 33096 28273 33099
rect 22152 33068 28273 33096
rect 22152 33056 22158 33068
rect 28261 33065 28273 33068
rect 28307 33065 28319 33099
rect 28261 33059 28319 33065
rect 18046 33028 18052 33040
rect 17788 33000 18052 33028
rect 17788 32969 17816 33000
rect 18046 32988 18052 33000
rect 18104 32988 18110 33040
rect 22738 33028 22744 33040
rect 22699 33000 22744 33028
rect 22738 32988 22744 33000
rect 22796 32988 22802 33040
rect 23290 33028 23296 33040
rect 23251 33000 23296 33028
rect 23290 32988 23296 33000
rect 23348 32988 23354 33040
rect 24394 33028 24400 33040
rect 24355 33000 24400 33028
rect 24394 32988 24400 33000
rect 24452 32988 24458 33040
rect 30469 33031 30527 33037
rect 30469 33028 30481 33031
rect 27908 33000 30481 33028
rect 17773 32963 17831 32969
rect 17773 32929 17785 32963
rect 17819 32929 17831 32963
rect 17773 32923 17831 32929
rect 17862 32920 17868 32972
rect 17920 32960 17926 32972
rect 17957 32963 18015 32969
rect 17957 32960 17969 32963
rect 17920 32932 17969 32960
rect 17920 32920 17926 32932
rect 17957 32929 17969 32932
rect 18003 32929 18015 32963
rect 17957 32923 18015 32929
rect 20070 32920 20076 32972
rect 20128 32960 20134 32972
rect 22094 32960 22100 32972
rect 20128 32932 22100 32960
rect 20128 32920 20134 32932
rect 22094 32920 22100 32932
rect 22152 32920 22158 32972
rect 22204 32932 23428 32960
rect 12710 32852 12716 32904
rect 12768 32892 12774 32904
rect 12805 32895 12863 32901
rect 12805 32892 12817 32895
rect 12768 32864 12817 32892
rect 12768 32852 12774 32864
rect 12805 32861 12817 32864
rect 12851 32861 12863 32895
rect 12805 32855 12863 32861
rect 12820 32824 12848 32855
rect 12894 32852 12900 32904
rect 12952 32892 12958 32904
rect 19242 32892 19248 32904
rect 12952 32864 19248 32892
rect 12952 32852 12958 32864
rect 19242 32852 19248 32864
rect 19300 32852 19306 32904
rect 22204 32892 22232 32932
rect 21284 32864 22232 32892
rect 23400 32892 23428 32932
rect 25700 32932 27016 32960
rect 25700 32892 25728 32932
rect 23400 32864 25728 32892
rect 13265 32827 13323 32833
rect 13265 32824 13277 32827
rect 12820 32796 13277 32824
rect 13265 32793 13277 32796
rect 13311 32793 13323 32827
rect 13265 32787 13323 32793
rect 18049 32827 18107 32833
rect 18049 32793 18061 32827
rect 18095 32824 18107 32827
rect 19150 32824 19156 32836
rect 18095 32796 19156 32824
rect 18095 32793 18107 32796
rect 18049 32787 18107 32793
rect 19150 32784 19156 32796
rect 19208 32824 19214 32836
rect 19337 32827 19395 32833
rect 19337 32824 19349 32827
rect 19208 32796 19349 32824
rect 19208 32784 19214 32796
rect 19337 32793 19349 32796
rect 19383 32824 19395 32827
rect 21284 32824 21312 32864
rect 25774 32852 25780 32904
rect 25832 32892 25838 32904
rect 26050 32892 26056 32904
rect 25832 32864 26056 32892
rect 25832 32852 25838 32864
rect 26050 32852 26056 32864
rect 26108 32892 26114 32904
rect 26881 32895 26939 32901
rect 26881 32892 26893 32895
rect 26108 32864 26893 32892
rect 26108 32852 26114 32864
rect 26881 32861 26893 32864
rect 26927 32861 26939 32895
rect 26988 32892 27016 32932
rect 27908 32892 27936 33000
rect 30469 32997 30481 33000
rect 30515 32997 30527 33031
rect 30469 32991 30527 32997
rect 26988 32864 27936 32892
rect 26881 32855 26939 32861
rect 28994 32852 29000 32904
rect 29052 32892 29058 32904
rect 31582 32895 31640 32901
rect 31582 32892 31594 32895
rect 29052 32864 31594 32892
rect 29052 32852 29058 32864
rect 31582 32861 31594 32864
rect 31628 32861 31640 32895
rect 31582 32855 31640 32861
rect 31849 32895 31907 32901
rect 31849 32861 31861 32895
rect 31895 32892 31907 32895
rect 33134 32892 33140 32904
rect 31895 32864 33140 32892
rect 31895 32861 31907 32864
rect 31849 32855 31907 32861
rect 33134 32852 33140 32864
rect 33192 32892 33198 32904
rect 33689 32895 33747 32901
rect 33689 32892 33701 32895
rect 33192 32864 33701 32892
rect 33192 32852 33198 32864
rect 33689 32861 33701 32864
rect 33735 32861 33747 32895
rect 33689 32855 33747 32861
rect 19383 32796 21312 32824
rect 19383 32793 19395 32796
rect 19337 32787 19395 32793
rect 21358 32784 21364 32836
rect 21416 32824 21422 32836
rect 24394 32824 24400 32836
rect 21416 32796 24400 32824
rect 21416 32784 21422 32796
rect 24394 32784 24400 32796
rect 24452 32784 24458 32836
rect 24486 32784 24492 32836
rect 24544 32824 24550 32836
rect 25510 32827 25568 32833
rect 25510 32824 25522 32827
rect 24544 32796 25522 32824
rect 24544 32784 24550 32796
rect 25510 32793 25522 32796
rect 25556 32793 25568 32827
rect 27126 32827 27184 32833
rect 27126 32824 27138 32827
rect 25510 32787 25568 32793
rect 25700 32796 27138 32824
rect 14182 32756 14188 32768
rect 14143 32728 14188 32756
rect 14182 32716 14188 32728
rect 14240 32716 14246 32768
rect 23106 32716 23112 32768
rect 23164 32756 23170 32768
rect 25700 32756 25728 32796
rect 27126 32793 27138 32796
rect 27172 32793 27184 32827
rect 27126 32787 27184 32793
rect 27246 32784 27252 32836
rect 27304 32824 27310 32836
rect 27304 32796 30604 32824
rect 27304 32784 27310 32796
rect 23164 32728 25728 32756
rect 30576 32756 30604 32796
rect 33318 32784 33324 32836
rect 33376 32824 33382 32836
rect 33422 32827 33480 32833
rect 33422 32824 33434 32827
rect 33376 32796 33434 32824
rect 33376 32784 33382 32796
rect 33422 32793 33434 32796
rect 33468 32793 33480 32827
rect 33422 32787 33480 32793
rect 32309 32759 32367 32765
rect 32309 32756 32321 32759
rect 30576 32728 32321 32756
rect 23164 32716 23170 32728
rect 32309 32725 32321 32728
rect 32355 32725 32367 32759
rect 32309 32719 32367 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 12437 32555 12495 32561
rect 12437 32521 12449 32555
rect 12483 32552 12495 32555
rect 12483 32524 23980 32552
rect 12483 32521 12495 32524
rect 12437 32515 12495 32521
rect 5074 32444 5080 32496
rect 5132 32484 5138 32496
rect 12894 32484 12900 32496
rect 5132 32456 12900 32484
rect 5132 32444 5138 32456
rect 12894 32444 12900 32456
rect 12952 32444 12958 32496
rect 13170 32484 13176 32496
rect 13131 32456 13176 32484
rect 13170 32444 13176 32456
rect 13228 32444 13234 32496
rect 14001 32487 14059 32493
rect 14001 32484 14013 32487
rect 13464 32456 14013 32484
rect 12250 32416 12256 32428
rect 12211 32388 12256 32416
rect 12250 32376 12256 32388
rect 12308 32376 12314 32428
rect 13464 32425 13492 32456
rect 14001 32453 14013 32456
rect 14047 32484 14059 32487
rect 14182 32484 14188 32496
rect 14047 32456 14188 32484
rect 14047 32453 14059 32456
rect 14001 32447 14059 32453
rect 14182 32444 14188 32456
rect 14240 32484 14246 32496
rect 14240 32456 14964 32484
rect 14240 32444 14246 32456
rect 13449 32419 13507 32425
rect 13449 32385 13461 32419
rect 13495 32385 13507 32419
rect 13906 32416 13912 32428
rect 13867 32388 13912 32416
rect 13449 32379 13507 32385
rect 13906 32376 13912 32388
rect 13964 32376 13970 32428
rect 14369 32419 14427 32425
rect 14369 32416 14381 32419
rect 14108 32388 14381 32416
rect 13173 32351 13231 32357
rect 13173 32317 13185 32351
rect 13219 32348 13231 32351
rect 14108 32348 14136 32388
rect 14369 32385 14381 32388
rect 14415 32385 14427 32419
rect 14369 32379 14427 32385
rect 14936 32357 14964 32456
rect 15010 32444 15016 32496
rect 15068 32484 15074 32496
rect 23382 32484 23388 32496
rect 15068 32456 23388 32484
rect 15068 32444 15074 32456
rect 23382 32444 23388 32456
rect 23440 32444 23446 32496
rect 23952 32484 23980 32524
rect 36262 32512 36268 32564
rect 36320 32552 36326 32564
rect 36357 32555 36415 32561
rect 36357 32552 36369 32555
rect 36320 32524 36369 32552
rect 36320 32512 36326 32524
rect 36357 32521 36369 32524
rect 36403 32521 36415 32555
rect 36357 32515 36415 32521
rect 25786 32487 25844 32493
rect 25786 32484 25798 32487
rect 23952 32456 25798 32484
rect 25786 32453 25798 32456
rect 25832 32453 25844 32487
rect 25786 32447 25844 32453
rect 25884 32456 31754 32484
rect 16758 32376 16764 32428
rect 16816 32416 16822 32428
rect 18233 32419 18291 32425
rect 18233 32416 18245 32419
rect 16816 32388 18245 32416
rect 16816 32376 16822 32388
rect 18233 32385 18245 32388
rect 18279 32416 18291 32419
rect 18969 32419 19027 32425
rect 18969 32416 18981 32419
rect 18279 32388 18981 32416
rect 18279 32385 18291 32388
rect 18233 32379 18291 32385
rect 18969 32385 18981 32388
rect 19015 32385 19027 32419
rect 18969 32379 19027 32385
rect 19153 32419 19211 32425
rect 19153 32385 19165 32419
rect 19199 32416 19211 32419
rect 19705 32419 19763 32425
rect 19705 32416 19717 32419
rect 19199 32388 19717 32416
rect 19199 32385 19211 32388
rect 19153 32379 19211 32385
rect 19705 32385 19717 32388
rect 19751 32385 19763 32419
rect 19705 32379 19763 32385
rect 22462 32376 22468 32428
rect 22520 32416 22526 32428
rect 22649 32419 22707 32425
rect 22649 32416 22661 32419
rect 22520 32388 22661 32416
rect 22520 32376 22526 32388
rect 22649 32385 22661 32388
rect 22695 32385 22707 32419
rect 25884 32416 25912 32456
rect 26050 32416 26056 32428
rect 22649 32379 22707 32385
rect 22848 32388 25912 32416
rect 26011 32388 26056 32416
rect 13219 32320 14136 32348
rect 14277 32351 14335 32357
rect 13219 32317 13231 32320
rect 13173 32311 13231 32317
rect 14277 32317 14289 32351
rect 14323 32317 14335 32351
rect 14277 32311 14335 32317
rect 14921 32351 14979 32357
rect 14921 32317 14933 32351
rect 14967 32348 14979 32351
rect 18782 32348 18788 32360
rect 14967 32320 18788 32348
rect 14967 32317 14979 32320
rect 14921 32311 14979 32317
rect 14292 32280 14320 32311
rect 18782 32308 18788 32320
rect 18840 32308 18846 32360
rect 16574 32280 16580 32292
rect 14292 32252 16580 32280
rect 16574 32240 16580 32252
rect 16632 32280 16638 32292
rect 17034 32280 17040 32292
rect 16632 32252 17040 32280
rect 16632 32240 16638 32252
rect 17034 32240 17040 32252
rect 17092 32240 17098 32292
rect 19889 32283 19947 32289
rect 19889 32249 19901 32283
rect 19935 32280 19947 32283
rect 22738 32280 22744 32292
rect 19935 32252 22744 32280
rect 19935 32249 19947 32252
rect 19889 32243 19947 32249
rect 22738 32240 22744 32252
rect 22796 32240 22802 32292
rect 22848 32289 22876 32388
rect 26050 32376 26056 32388
rect 26108 32376 26114 32428
rect 26142 32376 26148 32428
rect 26200 32416 26206 32428
rect 28914 32419 28972 32425
rect 28914 32416 28926 32419
rect 26200 32388 28926 32416
rect 26200 32376 26206 32388
rect 28914 32385 28926 32388
rect 28960 32385 28972 32419
rect 28914 32379 28972 32385
rect 29730 32376 29736 32428
rect 29788 32416 29794 32428
rect 29897 32419 29955 32425
rect 29897 32416 29909 32419
rect 29788 32388 29909 32416
rect 29788 32376 29794 32388
rect 29897 32385 29909 32388
rect 29943 32385 29955 32419
rect 31726 32416 31754 32456
rect 35233 32419 35291 32425
rect 35233 32416 35245 32419
rect 31726 32388 35245 32416
rect 29897 32379 29955 32385
rect 35233 32385 35245 32388
rect 35279 32385 35291 32419
rect 35233 32379 35291 32385
rect 29181 32351 29239 32357
rect 29181 32317 29193 32351
rect 29227 32348 29239 32351
rect 29638 32348 29644 32360
rect 29227 32320 29644 32348
rect 29227 32317 29239 32320
rect 29181 32311 29239 32317
rect 29638 32308 29644 32320
rect 29696 32308 29702 32360
rect 34977 32351 35035 32357
rect 34977 32317 34989 32351
rect 35023 32317 35035 32351
rect 34977 32311 35035 32317
rect 22833 32283 22891 32289
rect 22833 32249 22845 32283
rect 22879 32249 22891 32283
rect 31018 32280 31024 32292
rect 30979 32252 31024 32280
rect 22833 32243 22891 32249
rect 31018 32240 31024 32252
rect 31076 32240 31082 32292
rect 13357 32215 13415 32221
rect 13357 32181 13369 32215
rect 13403 32212 13415 32215
rect 13906 32212 13912 32224
rect 13403 32184 13912 32212
rect 13403 32181 13415 32184
rect 13357 32175 13415 32181
rect 13906 32172 13912 32184
rect 13964 32172 13970 32224
rect 14185 32215 14243 32221
rect 14185 32181 14197 32215
rect 14231 32212 14243 32215
rect 15930 32212 15936 32224
rect 14231 32184 15936 32212
rect 14231 32181 14243 32184
rect 14185 32175 14243 32181
rect 15930 32172 15936 32184
rect 15988 32212 15994 32224
rect 16482 32212 16488 32224
rect 15988 32184 16488 32212
rect 15988 32172 15994 32184
rect 16482 32172 16488 32184
rect 16540 32172 16546 32224
rect 21450 32172 21456 32224
rect 21508 32212 21514 32224
rect 21821 32215 21879 32221
rect 21821 32212 21833 32215
rect 21508 32184 21833 32212
rect 21508 32172 21514 32184
rect 21821 32181 21833 32184
rect 21867 32181 21879 32215
rect 24670 32212 24676 32224
rect 24631 32184 24676 32212
rect 21821 32175 21879 32181
rect 24670 32172 24676 32184
rect 24728 32172 24734 32224
rect 27614 32172 27620 32224
rect 27672 32212 27678 32224
rect 27801 32215 27859 32221
rect 27801 32212 27813 32215
rect 27672 32184 27813 32212
rect 27672 32172 27678 32184
rect 27801 32181 27813 32184
rect 27847 32181 27859 32215
rect 34992 32212 35020 32311
rect 35894 32212 35900 32224
rect 34992 32184 35900 32212
rect 27801 32175 27859 32181
rect 35894 32172 35900 32184
rect 35952 32172 35958 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 13541 32011 13599 32017
rect 13541 31977 13553 32011
rect 13587 32008 13599 32011
rect 13906 32008 13912 32020
rect 13587 31980 13912 32008
rect 13587 31977 13599 31980
rect 13541 31971 13599 31977
rect 13906 31968 13912 31980
rect 13964 32008 13970 32020
rect 14553 32011 14611 32017
rect 14553 32008 14565 32011
rect 13964 31980 14565 32008
rect 13964 31968 13970 31980
rect 14553 31977 14565 31980
rect 14599 32008 14611 32011
rect 15010 32008 15016 32020
rect 14599 31980 15016 32008
rect 14599 31977 14611 31980
rect 14553 31971 14611 31977
rect 15010 31968 15016 31980
rect 15068 31968 15074 32020
rect 16853 32011 16911 32017
rect 16853 31977 16865 32011
rect 16899 32008 16911 32011
rect 22189 32011 22247 32017
rect 16899 31980 21680 32008
rect 16899 31977 16911 31980
rect 16853 31971 16911 31977
rect 21358 31940 21364 31952
rect 15856 31912 21364 31940
rect 15856 31813 15884 31912
rect 21358 31900 21364 31912
rect 21416 31900 21422 31952
rect 21545 31943 21603 31949
rect 21545 31909 21557 31943
rect 21591 31909 21603 31943
rect 21652 31940 21680 31980
rect 22189 31977 22201 32011
rect 22235 32008 22247 32011
rect 26142 32008 26148 32020
rect 22235 31980 26148 32008
rect 22235 31977 22247 31980
rect 22189 31971 22247 31977
rect 26142 31968 26148 31980
rect 26200 31968 26206 32020
rect 29546 31968 29552 32020
rect 29604 32008 29610 32020
rect 29641 32011 29699 32017
rect 29641 32008 29653 32011
rect 29604 31980 29653 32008
rect 29604 31968 29610 31980
rect 29641 31977 29653 31980
rect 29687 32008 29699 32011
rect 29730 32008 29736 32020
rect 29687 31980 29736 32008
rect 29687 31977 29699 31980
rect 29641 31971 29699 31977
rect 29730 31968 29736 31980
rect 29788 31968 29794 32020
rect 31386 31968 31392 32020
rect 31444 32008 31450 32020
rect 34790 32008 34796 32020
rect 31444 31980 33272 32008
rect 34751 31980 34796 32008
rect 31444 31968 31450 31980
rect 24394 31940 24400 31952
rect 21652 31912 23796 31940
rect 24355 31912 24400 31940
rect 21545 31903 21603 31909
rect 15930 31832 15936 31884
rect 15988 31872 15994 31884
rect 16209 31875 16267 31881
rect 15988 31844 16033 31872
rect 15988 31832 15994 31844
rect 16209 31841 16221 31875
rect 16255 31872 16267 31875
rect 17126 31872 17132 31884
rect 16255 31844 17132 31872
rect 16255 31841 16267 31844
rect 16209 31835 16267 31841
rect 17126 31832 17132 31844
rect 17184 31832 17190 31884
rect 20714 31832 20720 31884
rect 20772 31872 20778 31884
rect 20901 31875 20959 31881
rect 20901 31872 20913 31875
rect 20772 31844 20913 31872
rect 20772 31832 20778 31844
rect 20901 31841 20913 31844
rect 20947 31841 20959 31875
rect 21082 31872 21088 31884
rect 21043 31844 21088 31872
rect 20901 31835 20959 31841
rect 21082 31832 21088 31844
rect 21140 31832 21146 31884
rect 21560 31872 21588 31903
rect 23768 31872 23796 31912
rect 24394 31900 24400 31912
rect 24452 31900 24458 31952
rect 31202 31900 31208 31952
rect 31260 31940 31266 31952
rect 31297 31943 31355 31949
rect 31297 31940 31309 31943
rect 31260 31912 31309 31940
rect 31260 31900 31266 31912
rect 31297 31909 31309 31912
rect 31343 31909 31355 31943
rect 31297 31903 31355 31909
rect 24762 31872 24768 31884
rect 21560 31844 22968 31872
rect 23768 31844 24768 31872
rect 15841 31807 15899 31813
rect 15841 31773 15853 31807
rect 15887 31773 15899 31807
rect 15841 31767 15899 31773
rect 16298 31764 16304 31816
rect 16356 31804 16362 31816
rect 16669 31807 16727 31813
rect 16669 31804 16681 31807
rect 16356 31776 16681 31804
rect 16356 31764 16362 31776
rect 16669 31773 16681 31776
rect 16715 31773 16727 31807
rect 16669 31767 16727 31773
rect 18782 31764 18788 31816
rect 18840 31804 18846 31816
rect 19337 31807 19395 31813
rect 19337 31804 19349 31807
rect 18840 31776 19349 31804
rect 18840 31764 18846 31776
rect 19337 31773 19349 31776
rect 19383 31804 19395 31807
rect 22002 31804 22008 31816
rect 19383 31776 21864 31804
rect 21963 31776 22008 31804
rect 19383 31773 19395 31776
rect 19337 31767 19395 31773
rect 21177 31739 21235 31745
rect 21177 31705 21189 31739
rect 21223 31736 21235 31739
rect 21450 31736 21456 31748
rect 21223 31708 21456 31736
rect 21223 31705 21235 31708
rect 21177 31699 21235 31705
rect 21450 31696 21456 31708
rect 21508 31696 21514 31748
rect 21836 31736 21864 31776
rect 22002 31764 22008 31776
rect 22060 31764 22066 31816
rect 22940 31813 22968 31844
rect 24762 31832 24768 31844
rect 24820 31832 24826 31884
rect 25777 31875 25835 31881
rect 25777 31841 25789 31875
rect 25823 31872 25835 31875
rect 26050 31872 26056 31884
rect 25823 31844 26056 31872
rect 25823 31841 25835 31844
rect 25777 31835 25835 31841
rect 26050 31832 26056 31844
rect 26108 31832 26114 31884
rect 22925 31807 22983 31813
rect 22112 31776 22784 31804
rect 22112 31736 22140 31776
rect 21836 31708 22140 31736
rect 22756 31736 22784 31776
rect 22925 31773 22937 31807
rect 22971 31773 22983 31807
rect 24946 31804 24952 31816
rect 22925 31767 22983 31773
rect 23032 31776 24952 31804
rect 23032 31736 23060 31776
rect 24946 31764 24952 31776
rect 25004 31764 25010 31816
rect 25038 31764 25044 31816
rect 25096 31804 25102 31816
rect 25510 31807 25568 31813
rect 25510 31804 25522 31807
rect 25096 31776 25522 31804
rect 25096 31764 25102 31776
rect 25510 31773 25522 31776
rect 25556 31773 25568 31807
rect 25510 31767 25568 31773
rect 32677 31807 32735 31813
rect 32677 31773 32689 31807
rect 32723 31804 32735 31807
rect 33134 31804 33140 31816
rect 32723 31776 33140 31804
rect 32723 31773 32735 31776
rect 32677 31767 32735 31773
rect 33134 31764 33140 31776
rect 33192 31764 33198 31816
rect 33244 31804 33272 31980
rect 34790 31968 34796 31980
rect 34848 31968 34854 32020
rect 38105 32011 38163 32017
rect 38105 32008 38117 32011
rect 35866 31980 38117 32008
rect 34698 31900 34704 31952
rect 34756 31940 34762 31952
rect 35866 31940 35894 31980
rect 38105 31977 38117 31980
rect 38151 31977 38163 32011
rect 38105 31971 38163 31977
rect 34756 31912 35894 31940
rect 34756 31900 34762 31912
rect 35894 31832 35900 31884
rect 35952 31872 35958 31884
rect 36725 31875 36783 31881
rect 36725 31872 36737 31875
rect 35952 31844 36737 31872
rect 35952 31832 35958 31844
rect 36725 31841 36737 31844
rect 36771 31841 36783 31875
rect 36725 31835 36783 31841
rect 36981 31807 37039 31813
rect 36981 31804 36993 31807
rect 33244 31776 36993 31804
rect 36981 31773 36993 31776
rect 37027 31773 37039 31807
rect 36981 31767 37039 31773
rect 22756 31708 23060 31736
rect 32410 31739 32468 31745
rect 32410 31705 32422 31739
rect 32456 31705 32468 31739
rect 32410 31699 32468 31705
rect 23106 31668 23112 31680
rect 23067 31640 23112 31668
rect 23106 31628 23112 31640
rect 23164 31628 23170 31680
rect 30650 31628 30656 31680
rect 30708 31668 30714 31680
rect 30745 31671 30803 31677
rect 30745 31668 30757 31671
rect 30708 31640 30757 31668
rect 30708 31628 30714 31640
rect 30745 31637 30757 31640
rect 30791 31668 30803 31671
rect 32425 31668 32453 31699
rect 35250 31668 35256 31680
rect 30791 31640 32453 31668
rect 35211 31640 35256 31668
rect 30791 31637 30803 31640
rect 30745 31631 30803 31637
rect 35250 31628 35256 31640
rect 35308 31628 35314 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 27614 31464 27620 31476
rect 18708 31436 27620 31464
rect 16666 31328 16672 31340
rect 16627 31300 16672 31328
rect 16666 31288 16672 31300
rect 16724 31288 16730 31340
rect 18708 31337 18736 31436
rect 27614 31424 27620 31436
rect 27672 31424 27678 31476
rect 34882 31424 34888 31476
rect 34940 31464 34946 31476
rect 35618 31464 35624 31476
rect 34940 31436 35624 31464
rect 34940 31424 34946 31436
rect 35618 31424 35624 31436
rect 35676 31424 35682 31476
rect 20346 31356 20352 31408
rect 20404 31396 20410 31408
rect 22097 31399 22155 31405
rect 22097 31396 22109 31399
rect 20404 31368 22109 31396
rect 20404 31356 20410 31368
rect 22097 31365 22109 31368
rect 22143 31365 22155 31399
rect 22097 31359 22155 31365
rect 23106 31356 23112 31408
rect 23164 31396 23170 31408
rect 25418 31399 25476 31405
rect 25418 31396 25430 31399
rect 23164 31368 25430 31396
rect 23164 31356 23170 31368
rect 25418 31365 25430 31368
rect 25464 31365 25476 31399
rect 25418 31359 25476 31365
rect 25590 31356 25596 31408
rect 25648 31396 25654 31408
rect 27218 31399 27276 31405
rect 27218 31396 27230 31399
rect 25648 31368 27230 31396
rect 25648 31356 25654 31368
rect 27218 31365 27230 31368
rect 27264 31365 27276 31399
rect 27218 31359 27276 31365
rect 29638 31356 29644 31408
rect 29696 31396 29702 31408
rect 34241 31399 34299 31405
rect 29696 31368 30512 31396
rect 29696 31356 29702 31368
rect 18693 31331 18751 31337
rect 18693 31297 18705 31331
rect 18739 31297 18751 31331
rect 20438 31328 20444 31340
rect 20399 31300 20444 31328
rect 18693 31291 18751 31297
rect 20438 31288 20444 31300
rect 20496 31288 20502 31340
rect 22189 31331 22247 31337
rect 22189 31297 22201 31331
rect 22235 31328 22247 31331
rect 23017 31331 23075 31337
rect 23017 31328 23029 31331
rect 22235 31300 23029 31328
rect 22235 31297 22247 31300
rect 22189 31291 22247 31297
rect 23017 31297 23029 31300
rect 23063 31328 23075 31331
rect 24394 31328 24400 31340
rect 23063 31300 24400 31328
rect 23063 31297 23075 31300
rect 23017 31291 23075 31297
rect 24394 31288 24400 31300
rect 24452 31288 24458 31340
rect 25685 31331 25743 31337
rect 25685 31297 25697 31331
rect 25731 31328 25743 31331
rect 26050 31328 26056 31340
rect 25731 31300 26056 31328
rect 25731 31297 25743 31300
rect 25685 31291 25743 31297
rect 26050 31288 26056 31300
rect 26108 31328 26114 31340
rect 26973 31331 27031 31337
rect 26973 31328 26985 31331
rect 26108 31300 26985 31328
rect 26108 31288 26114 31300
rect 26973 31297 26985 31300
rect 27019 31297 27031 31331
rect 26973 31291 27031 31297
rect 28994 31288 29000 31340
rect 29052 31328 29058 31340
rect 30484 31337 30512 31368
rect 34241 31365 34253 31399
rect 34287 31396 34299 31399
rect 34790 31396 34796 31408
rect 34287 31368 34796 31396
rect 34287 31365 34299 31368
rect 34241 31359 34299 31365
rect 34790 31356 34796 31368
rect 34848 31356 34854 31408
rect 30202 31331 30260 31337
rect 30202 31328 30214 31331
rect 29052 31300 30214 31328
rect 29052 31288 29058 31300
rect 30202 31297 30214 31300
rect 30248 31297 30260 31331
rect 30202 31291 30260 31297
rect 30469 31331 30527 31337
rect 30469 31297 30481 31331
rect 30515 31297 30527 31331
rect 30469 31291 30527 31297
rect 33134 31288 33140 31340
rect 33192 31328 33198 31340
rect 34701 31331 34759 31337
rect 34701 31328 34713 31331
rect 33192 31300 34713 31328
rect 33192 31288 33198 31300
rect 34701 31297 34713 31300
rect 34747 31297 34759 31331
rect 34957 31331 35015 31337
rect 34957 31328 34969 31331
rect 34701 31291 34759 31297
rect 34808 31300 34969 31328
rect 17034 31220 17040 31272
rect 17092 31260 17098 31272
rect 18601 31263 18659 31269
rect 18601 31260 18613 31263
rect 17092 31232 18613 31260
rect 17092 31220 17098 31232
rect 18601 31229 18613 31232
rect 18647 31229 18659 31263
rect 18601 31223 18659 31229
rect 19061 31263 19119 31269
rect 19061 31229 19073 31263
rect 19107 31260 19119 31263
rect 20714 31260 20720 31272
rect 19107 31232 20720 31260
rect 19107 31229 19119 31232
rect 19061 31223 19119 31229
rect 20714 31220 20720 31232
rect 20772 31220 20778 31272
rect 20806 31220 20812 31272
rect 20864 31260 20870 31272
rect 21910 31260 21916 31272
rect 20864 31232 21916 31260
rect 20864 31220 20870 31232
rect 21910 31220 21916 31232
rect 21968 31220 21974 31272
rect 22066 31232 24624 31260
rect 4706 31152 4712 31204
rect 4764 31192 4770 31204
rect 16853 31195 16911 31201
rect 4764 31164 6914 31192
rect 4764 31152 4770 31164
rect 6886 31124 6914 31164
rect 16853 31161 16865 31195
rect 16899 31192 16911 31195
rect 22066 31192 22094 31232
rect 24486 31192 24492 31204
rect 16899 31164 22094 31192
rect 22388 31164 24492 31192
rect 16899 31161 16911 31164
rect 16853 31155 16911 31161
rect 17770 31124 17776 31136
rect 6886 31096 17776 31124
rect 17770 31084 17776 31096
rect 17828 31084 17834 31136
rect 17954 31124 17960 31136
rect 17915 31096 17960 31124
rect 17954 31084 17960 31096
rect 18012 31124 18018 31136
rect 18138 31124 18144 31136
rect 18012 31096 18144 31124
rect 18012 31084 18018 31096
rect 18138 31084 18144 31096
rect 18196 31084 18202 31136
rect 20625 31127 20683 31133
rect 20625 31093 20637 31127
rect 20671 31124 20683 31127
rect 22388 31124 22416 31164
rect 24486 31152 24492 31164
rect 24544 31152 24550 31204
rect 24596 31192 24624 31232
rect 34606 31220 34612 31272
rect 34664 31260 34670 31272
rect 34808 31260 34836 31300
rect 34957 31297 34969 31300
rect 35003 31328 35015 31331
rect 35250 31328 35256 31340
rect 35003 31300 35256 31328
rect 35003 31297 35015 31300
rect 34957 31291 35015 31297
rect 35250 31288 35256 31300
rect 35308 31288 35314 31340
rect 34664 31232 34836 31260
rect 34664 31220 34670 31232
rect 24596 31164 24808 31192
rect 22554 31124 22560 31136
rect 20671 31096 22416 31124
rect 22515 31096 22560 31124
rect 20671 31093 20683 31096
rect 20625 31087 20683 31093
rect 22554 31084 22560 31096
rect 22612 31084 22618 31136
rect 24302 31124 24308 31136
rect 24263 31096 24308 31124
rect 24302 31084 24308 31096
rect 24360 31084 24366 31136
rect 24780 31124 24808 31164
rect 28074 31124 28080 31136
rect 24780 31096 28080 31124
rect 28074 31084 28080 31096
rect 28132 31084 28138 31136
rect 28350 31124 28356 31136
rect 28311 31096 28356 31124
rect 28350 31084 28356 31096
rect 28408 31084 28414 31136
rect 29086 31124 29092 31136
rect 29047 31096 29092 31124
rect 29086 31084 29092 31096
rect 29144 31084 29150 31136
rect 32953 31127 33011 31133
rect 32953 31093 32965 31127
rect 32999 31124 33011 31127
rect 33134 31124 33140 31136
rect 32999 31096 33140 31124
rect 32999 31093 33011 31096
rect 32953 31087 33011 31093
rect 33134 31084 33140 31096
rect 33192 31084 33198 31136
rect 36078 31124 36084 31136
rect 36039 31096 36084 31124
rect 36078 31084 36084 31096
rect 36136 31084 36142 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 12161 30923 12219 30929
rect 12161 30889 12173 30923
rect 12207 30920 12219 30923
rect 12250 30920 12256 30932
rect 12207 30892 12256 30920
rect 12207 30889 12219 30892
rect 12161 30883 12219 30889
rect 12250 30880 12256 30892
rect 12308 30880 12314 30932
rect 17770 30880 17776 30932
rect 17828 30920 17834 30932
rect 18417 30923 18475 30929
rect 17828 30892 18368 30920
rect 17828 30880 17834 30892
rect 18046 30852 18052 30864
rect 17052 30824 18052 30852
rect 17052 30793 17080 30824
rect 18046 30812 18052 30824
rect 18104 30812 18110 30864
rect 18340 30852 18368 30892
rect 18417 30889 18429 30923
rect 18463 30920 18475 30923
rect 20438 30920 20444 30932
rect 18463 30892 20444 30920
rect 18463 30889 18475 30892
rect 18417 30883 18475 30889
rect 20438 30880 20444 30892
rect 20496 30880 20502 30932
rect 20901 30923 20959 30929
rect 20901 30889 20913 30923
rect 20947 30920 20959 30923
rect 22002 30920 22008 30932
rect 20947 30892 22008 30920
rect 20947 30889 20959 30892
rect 20901 30883 20959 30889
rect 22002 30880 22008 30892
rect 22060 30880 22066 30932
rect 30929 30923 30987 30929
rect 30929 30889 30941 30923
rect 30975 30920 30987 30923
rect 32122 30920 32128 30932
rect 30975 30892 32128 30920
rect 30975 30889 30987 30892
rect 30929 30883 30987 30889
rect 32122 30880 32128 30892
rect 32180 30880 32186 30932
rect 36446 30920 36452 30932
rect 36407 30892 36452 30920
rect 36446 30880 36452 30892
rect 36504 30880 36510 30932
rect 19978 30852 19984 30864
rect 18340 30824 19984 30852
rect 19978 30812 19984 30824
rect 20036 30812 20042 30864
rect 21542 30812 21548 30864
rect 21600 30852 21606 30864
rect 24302 30852 24308 30864
rect 21600 30824 24308 30852
rect 21600 30812 21606 30824
rect 24302 30812 24308 30824
rect 24360 30812 24366 30864
rect 17037 30787 17095 30793
rect 17037 30753 17049 30787
rect 17083 30753 17095 30787
rect 17037 30747 17095 30753
rect 17126 30744 17132 30796
rect 17184 30784 17190 30796
rect 26050 30784 26056 30796
rect 17184 30756 18276 30784
rect 26011 30756 26056 30784
rect 17184 30744 17190 30756
rect 11790 30716 11796 30728
rect 11751 30688 11796 30716
rect 11790 30676 11796 30688
rect 11848 30676 11854 30728
rect 11974 30716 11980 30728
rect 11935 30688 11980 30716
rect 11974 30676 11980 30688
rect 12032 30676 12038 30728
rect 12618 30716 12624 30728
rect 12579 30688 12624 30716
rect 12618 30676 12624 30688
rect 12676 30676 12682 30728
rect 17954 30676 17960 30728
rect 18012 30716 18018 30728
rect 18248 30725 18276 30756
rect 26050 30744 26056 30756
rect 26108 30744 26114 30796
rect 18141 30719 18199 30725
rect 18141 30716 18153 30719
rect 18012 30688 18153 30716
rect 18012 30676 18018 30688
rect 18141 30685 18153 30688
rect 18187 30685 18199 30719
rect 18141 30679 18199 30685
rect 18233 30719 18291 30725
rect 18233 30685 18245 30719
rect 18279 30685 18291 30719
rect 18233 30679 18291 30685
rect 20073 30719 20131 30725
rect 20073 30685 20085 30719
rect 20119 30716 20131 30719
rect 20530 30716 20536 30728
rect 20119 30688 20536 30716
rect 20119 30685 20131 30688
rect 20073 30679 20131 30685
rect 17221 30651 17279 30657
rect 17221 30617 17233 30651
rect 17267 30648 17279 30651
rect 18046 30648 18052 30660
rect 17267 30620 18052 30648
rect 17267 30617 17279 30620
rect 17221 30611 17279 30617
rect 18046 30608 18052 30620
rect 18104 30608 18110 30660
rect 18156 30648 18184 30679
rect 20088 30648 20116 30679
rect 20530 30676 20536 30688
rect 20588 30676 20594 30728
rect 20714 30716 20720 30728
rect 20675 30688 20720 30716
rect 20714 30676 20720 30688
rect 20772 30676 20778 30728
rect 27798 30716 27804 30728
rect 27759 30688 27804 30716
rect 27798 30676 27804 30688
rect 27856 30676 27862 30728
rect 32306 30716 32312 30728
rect 32267 30688 32312 30716
rect 32306 30676 32312 30688
rect 32364 30676 32370 30728
rect 35069 30719 35127 30725
rect 35069 30685 35081 30719
rect 35115 30716 35127 30719
rect 35894 30716 35900 30728
rect 35115 30688 35900 30716
rect 35115 30685 35127 30688
rect 35069 30679 35127 30685
rect 35894 30676 35900 30688
rect 35952 30676 35958 30728
rect 18156 30620 20116 30648
rect 32042 30651 32100 30657
rect 32042 30617 32054 30651
rect 32088 30617 32100 30651
rect 32042 30611 32100 30617
rect 35336 30651 35394 30657
rect 35336 30617 35348 30651
rect 35382 30648 35394 30651
rect 35710 30648 35716 30660
rect 35382 30620 35716 30648
rect 35382 30617 35394 30620
rect 35336 30611 35394 30617
rect 12802 30580 12808 30592
rect 12763 30552 12808 30580
rect 12802 30540 12808 30552
rect 12860 30540 12866 30592
rect 17586 30580 17592 30592
rect 17547 30552 17592 30580
rect 17586 30540 17592 30552
rect 17644 30540 17650 30592
rect 32048 30580 32076 30611
rect 35710 30608 35716 30620
rect 35768 30608 35774 30660
rect 32122 30580 32128 30592
rect 32048 30552 32128 30580
rect 32122 30540 32128 30552
rect 32180 30540 32186 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 12802 30336 12808 30388
rect 12860 30376 12866 30388
rect 12860 30348 25553 30376
rect 12860 30336 12866 30348
rect 11885 30311 11943 30317
rect 11885 30277 11897 30311
rect 11931 30308 11943 30311
rect 12618 30308 12624 30320
rect 11931 30280 12624 30308
rect 11931 30277 11943 30280
rect 11885 30271 11943 30277
rect 12618 30268 12624 30280
rect 12676 30268 12682 30320
rect 15473 30311 15531 30317
rect 15473 30277 15485 30311
rect 15519 30308 15531 30311
rect 16666 30308 16672 30320
rect 15519 30280 16672 30308
rect 15519 30277 15531 30280
rect 15473 30271 15531 30277
rect 16666 30268 16672 30280
rect 16724 30268 16730 30320
rect 20530 30268 20536 30320
rect 20588 30308 20594 30320
rect 22186 30308 22192 30320
rect 20588 30280 22192 30308
rect 20588 30268 20594 30280
rect 22186 30268 22192 30280
rect 22244 30308 22250 30320
rect 25525 30317 25553 30348
rect 22373 30311 22431 30317
rect 22373 30308 22385 30311
rect 22244 30280 22385 30308
rect 22244 30268 22250 30280
rect 22373 30277 22385 30280
rect 22419 30277 22431 30311
rect 22373 30271 22431 30277
rect 25510 30311 25568 30317
rect 25510 30277 25522 30311
rect 25556 30277 25568 30311
rect 28994 30308 29000 30320
rect 25510 30271 25568 30277
rect 26160 30280 29000 30308
rect 11701 30243 11759 30249
rect 11701 30209 11713 30243
rect 11747 30240 11759 30243
rect 12250 30240 12256 30252
rect 11747 30212 12256 30240
rect 11747 30209 11759 30212
rect 11701 30203 11759 30209
rect 12250 30200 12256 30212
rect 12308 30200 12314 30252
rect 13725 30243 13783 30249
rect 13725 30209 13737 30243
rect 13771 30240 13783 30243
rect 14366 30240 14372 30252
rect 13771 30212 14372 30240
rect 13771 30209 13783 30212
rect 13725 30203 13783 30209
rect 14366 30200 14372 30212
rect 14424 30240 14430 30252
rect 15010 30240 15016 30252
rect 14424 30212 15016 30240
rect 14424 30200 14430 30212
rect 15010 30200 15016 30212
rect 15068 30200 15074 30252
rect 15286 30240 15292 30252
rect 15247 30212 15292 30240
rect 15286 30200 15292 30212
rect 15344 30200 15350 30252
rect 17494 30240 17500 30252
rect 17455 30212 17500 30240
rect 17494 30200 17500 30212
rect 17552 30200 17558 30252
rect 21726 30200 21732 30252
rect 21784 30240 21790 30252
rect 26160 30240 26188 30280
rect 28994 30268 29000 30280
rect 29052 30268 29058 30320
rect 21784 30212 26188 30240
rect 21784 30200 21790 30212
rect 27614 30200 27620 30252
rect 27672 30240 27678 30252
rect 28178 30243 28236 30249
rect 28178 30240 28190 30243
rect 27672 30212 28190 30240
rect 27672 30200 27678 30212
rect 28178 30209 28190 30212
rect 28224 30209 28236 30243
rect 28178 30203 28236 30209
rect 28350 30200 28356 30252
rect 28408 30240 28414 30252
rect 29161 30243 29219 30249
rect 29161 30240 29173 30243
rect 28408 30212 29173 30240
rect 28408 30200 28414 30212
rect 29161 30209 29173 30212
rect 29207 30209 29219 30243
rect 29161 30203 29219 30209
rect 33410 30200 33416 30252
rect 33468 30240 33474 30252
rect 34618 30243 34676 30249
rect 34618 30240 34630 30243
rect 33468 30212 34630 30240
rect 33468 30200 33474 30212
rect 34618 30209 34630 30212
rect 34664 30209 34676 30243
rect 34618 30203 34676 30209
rect 11517 30175 11575 30181
rect 11517 30141 11529 30175
rect 11563 30172 11575 30175
rect 11790 30172 11796 30184
rect 11563 30144 11796 30172
rect 11563 30141 11575 30144
rect 11517 30135 11575 30141
rect 11790 30132 11796 30144
rect 11848 30172 11854 30184
rect 15105 30175 15163 30181
rect 11848 30144 14320 30172
rect 11848 30132 11854 30144
rect 12618 29996 12624 30048
rect 12676 30036 12682 30048
rect 14292 30045 14320 30144
rect 15105 30141 15117 30175
rect 15151 30172 15163 30175
rect 15194 30172 15200 30184
rect 15151 30144 15200 30172
rect 15151 30141 15163 30144
rect 15105 30135 15163 30141
rect 15194 30132 15200 30144
rect 15252 30132 15258 30184
rect 25777 30175 25835 30181
rect 25777 30141 25789 30175
rect 25823 30172 25835 30175
rect 26510 30172 26516 30184
rect 25823 30144 26516 30172
rect 25823 30141 25835 30144
rect 25777 30135 25835 30141
rect 26510 30132 26516 30144
rect 26568 30132 26574 30184
rect 28445 30175 28503 30181
rect 28445 30141 28457 30175
rect 28491 30172 28503 30175
rect 28905 30175 28963 30181
rect 28905 30172 28917 30175
rect 28491 30144 28917 30172
rect 28491 30141 28503 30144
rect 28445 30135 28503 30141
rect 28905 30141 28917 30144
rect 28951 30141 28963 30175
rect 28905 30135 28963 30141
rect 34885 30175 34943 30181
rect 34885 30141 34897 30175
rect 34931 30172 34943 30175
rect 35894 30172 35900 30184
rect 34931 30144 35900 30172
rect 34931 30141 34943 30144
rect 34885 30135 34943 30141
rect 17681 30107 17739 30113
rect 17681 30073 17693 30107
rect 17727 30104 17739 30107
rect 17727 30076 24716 30104
rect 17727 30073 17739 30076
rect 17681 30067 17739 30073
rect 13081 30039 13139 30045
rect 13081 30036 13093 30039
rect 12676 30008 13093 30036
rect 12676 29996 12682 30008
rect 13081 30005 13093 30008
rect 13127 30005 13139 30039
rect 13081 29999 13139 30005
rect 14277 30039 14335 30045
rect 14277 30005 14289 30039
rect 14323 30036 14335 30039
rect 14366 30036 14372 30048
rect 14323 30008 14372 30036
rect 14323 30005 14335 30008
rect 14277 29999 14335 30005
rect 14366 29996 14372 30008
rect 14424 29996 14430 30048
rect 18046 29996 18052 30048
rect 18104 30036 18110 30048
rect 18233 30039 18291 30045
rect 18233 30036 18245 30039
rect 18104 30008 18245 30036
rect 18104 29996 18110 30008
rect 18233 30005 18245 30008
rect 18279 30036 18291 30039
rect 18598 30036 18604 30048
rect 18279 30008 18604 30036
rect 18279 30005 18291 30008
rect 18233 29999 18291 30005
rect 18598 29996 18604 30008
rect 18656 29996 18662 30048
rect 21913 30039 21971 30045
rect 21913 30005 21925 30039
rect 21959 30036 21971 30039
rect 22094 30036 22100 30048
rect 21959 30008 22100 30036
rect 21959 30005 21971 30008
rect 21913 29999 21971 30005
rect 22094 29996 22100 30008
rect 22152 29996 22158 30048
rect 24394 30036 24400 30048
rect 24355 30008 24400 30036
rect 24394 29996 24400 30008
rect 24452 29996 24458 30048
rect 24688 30036 24716 30076
rect 25866 30064 25872 30116
rect 25924 30104 25930 30116
rect 26326 30104 26332 30116
rect 25924 30076 26332 30104
rect 25924 30064 25930 30076
rect 26326 30064 26332 30076
rect 26384 30064 26390 30116
rect 25590 30036 25596 30048
rect 24688 30008 25596 30036
rect 25590 29996 25596 30008
rect 25648 29996 25654 30048
rect 26418 29996 26424 30048
rect 26476 30036 26482 30048
rect 27065 30039 27123 30045
rect 27065 30036 27077 30039
rect 26476 30008 27077 30036
rect 26476 29996 26482 30008
rect 27065 30005 27077 30008
rect 27111 30005 27123 30039
rect 28920 30036 28948 30135
rect 35894 30132 35900 30144
rect 35952 30132 35958 30184
rect 29270 30036 29276 30048
rect 28920 30008 29276 30036
rect 27065 29999 27123 30005
rect 29270 29996 29276 30008
rect 29328 29996 29334 30048
rect 30282 30036 30288 30048
rect 30243 30008 30288 30036
rect 30282 29996 30288 30008
rect 30340 29996 30346 30048
rect 33502 30036 33508 30048
rect 33463 30008 33508 30036
rect 33502 29996 33508 30008
rect 33560 29996 33566 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 11974 29792 11980 29844
rect 12032 29832 12038 29844
rect 12253 29835 12311 29841
rect 12253 29832 12265 29835
rect 12032 29804 12265 29832
rect 12032 29792 12038 29804
rect 12253 29801 12265 29804
rect 12299 29801 12311 29835
rect 16482 29832 16488 29844
rect 16443 29804 16488 29832
rect 12253 29795 12311 29801
rect 16482 29792 16488 29804
rect 16540 29792 16546 29844
rect 24394 29832 24400 29844
rect 16592 29804 24400 29832
rect 13538 29764 13544 29776
rect 13499 29736 13544 29764
rect 13538 29724 13544 29736
rect 13596 29724 13602 29776
rect 13722 29724 13728 29776
rect 13780 29764 13786 29776
rect 16592 29764 16620 29804
rect 24394 29792 24400 29804
rect 24452 29792 24458 29844
rect 25130 29792 25136 29844
rect 25188 29832 25194 29844
rect 25958 29832 25964 29844
rect 25188 29804 25964 29832
rect 25188 29792 25194 29804
rect 25958 29792 25964 29804
rect 26016 29832 26022 29844
rect 30282 29832 30288 29844
rect 26016 29804 30288 29832
rect 26016 29792 26022 29804
rect 30282 29792 30288 29804
rect 30340 29792 30346 29844
rect 33502 29832 33508 29844
rect 30392 29804 33508 29832
rect 22002 29764 22008 29776
rect 13780 29736 16620 29764
rect 21192 29736 22008 29764
rect 13780 29724 13786 29736
rect 12802 29696 12808 29708
rect 12763 29668 12808 29696
rect 12802 29656 12808 29668
rect 12860 29696 12866 29708
rect 15749 29699 15807 29705
rect 15749 29696 15761 29699
rect 12860 29668 15761 29696
rect 12860 29656 12866 29668
rect 15749 29665 15761 29668
rect 15795 29696 15807 29699
rect 15930 29696 15936 29708
rect 15795 29668 15936 29696
rect 15795 29665 15807 29668
rect 15749 29659 15807 29665
rect 15930 29656 15936 29668
rect 15988 29656 15994 29708
rect 21192 29696 21220 29736
rect 22002 29724 22008 29736
rect 22060 29724 22066 29776
rect 28902 29724 28908 29776
rect 28960 29764 28966 29776
rect 30392 29764 30420 29804
rect 33502 29792 33508 29804
rect 33560 29792 33566 29844
rect 36170 29792 36176 29844
rect 36228 29832 36234 29844
rect 36265 29835 36323 29841
rect 36265 29832 36277 29835
rect 36228 29804 36277 29832
rect 36228 29792 36234 29804
rect 36265 29801 36277 29804
rect 36311 29801 36323 29835
rect 36265 29795 36323 29801
rect 37918 29792 37924 29844
rect 37976 29832 37982 29844
rect 38102 29832 38108 29844
rect 37976 29804 38108 29832
rect 37976 29792 37982 29804
rect 38102 29792 38108 29804
rect 38160 29792 38166 29844
rect 28960 29736 30420 29764
rect 28960 29724 28966 29736
rect 21100 29668 21220 29696
rect 21288 29699 21346 29705
rect 21100 29640 21128 29668
rect 21288 29665 21300 29699
rect 21334 29696 21346 29699
rect 21726 29696 21732 29708
rect 21334 29668 21732 29696
rect 21334 29665 21346 29668
rect 21288 29659 21346 29665
rect 21726 29656 21732 29668
rect 21784 29656 21790 29708
rect 21821 29699 21879 29705
rect 21821 29665 21833 29699
rect 21867 29696 21879 29699
rect 22186 29696 22192 29708
rect 21867 29668 22192 29696
rect 21867 29665 21879 29668
rect 21821 29659 21879 29665
rect 22186 29656 22192 29668
rect 22244 29656 22250 29708
rect 32033 29699 32091 29705
rect 22388 29668 23336 29696
rect 12618 29588 12624 29640
rect 12676 29628 12682 29640
rect 12713 29631 12771 29637
rect 12713 29628 12725 29631
rect 12676 29600 12725 29628
rect 12676 29588 12682 29600
rect 12713 29597 12725 29600
rect 12759 29597 12771 29631
rect 14090 29628 14096 29640
rect 14051 29600 14096 29628
rect 12713 29591 12771 29597
rect 14090 29588 14096 29600
rect 14148 29588 14154 29640
rect 15565 29631 15623 29637
rect 15565 29597 15577 29631
rect 15611 29628 15623 29631
rect 16482 29628 16488 29640
rect 15611 29600 16488 29628
rect 15611 29597 15623 29600
rect 15565 29591 15623 29597
rect 16482 29588 16488 29600
rect 16540 29588 16546 29640
rect 17037 29631 17095 29637
rect 17037 29597 17049 29631
rect 17083 29628 17095 29631
rect 17586 29628 17592 29640
rect 17083 29600 17592 29628
rect 17083 29597 17095 29600
rect 17037 29591 17095 29597
rect 17586 29588 17592 29600
rect 17644 29588 17650 29640
rect 21082 29628 21088 29640
rect 20995 29600 21088 29628
rect 21082 29588 21088 29600
rect 21140 29588 21146 29640
rect 22094 29588 22100 29640
rect 22152 29628 22158 29640
rect 22388 29628 22416 29668
rect 22554 29628 22560 29640
rect 22152 29600 22416 29628
rect 22515 29600 22560 29628
rect 22152 29588 22158 29600
rect 22554 29588 22560 29600
rect 22612 29588 22618 29640
rect 23308 29637 23336 29668
rect 32033 29665 32045 29699
rect 32079 29696 32091 29699
rect 32306 29696 32312 29708
rect 32079 29668 32312 29696
rect 32079 29665 32091 29668
rect 32033 29659 32091 29665
rect 32306 29656 32312 29668
rect 32364 29656 32370 29708
rect 23293 29631 23351 29637
rect 23293 29597 23305 29631
rect 23339 29628 23351 29631
rect 25777 29631 25835 29637
rect 23339 29600 25636 29628
rect 23339 29597 23351 29600
rect 23293 29591 23351 29597
rect 10134 29520 10140 29572
rect 10192 29560 10198 29572
rect 20990 29560 20996 29572
rect 10192 29532 20996 29560
rect 10192 29520 10198 29532
rect 20990 29520 20996 29532
rect 21048 29520 21054 29572
rect 21361 29563 21419 29569
rect 21361 29529 21373 29563
rect 21407 29560 21419 29563
rect 21821 29563 21879 29569
rect 21821 29560 21833 29563
rect 21407 29532 21833 29560
rect 21407 29529 21419 29532
rect 21361 29523 21419 29529
rect 21821 29529 21833 29532
rect 21867 29529 21879 29563
rect 21821 29523 21879 29529
rect 24854 29520 24860 29572
rect 24912 29560 24918 29572
rect 25510 29563 25568 29569
rect 25510 29560 25522 29563
rect 24912 29532 25522 29560
rect 24912 29520 24918 29532
rect 25510 29529 25522 29532
rect 25556 29529 25568 29563
rect 25608 29560 25636 29600
rect 25777 29597 25789 29631
rect 25823 29628 25835 29631
rect 26510 29628 26516 29640
rect 25823 29600 26516 29628
rect 25823 29597 25835 29600
rect 25777 29591 25835 29597
rect 26510 29588 26516 29600
rect 26568 29588 26574 29640
rect 34885 29631 34943 29637
rect 34885 29597 34897 29631
rect 34931 29628 34943 29631
rect 35894 29628 35900 29640
rect 34931 29600 35900 29628
rect 34931 29597 34943 29600
rect 34885 29591 34943 29597
rect 35894 29588 35900 29600
rect 35952 29628 35958 29640
rect 36725 29631 36783 29637
rect 36725 29628 36737 29631
rect 35952 29600 36737 29628
rect 35952 29588 35958 29600
rect 36725 29597 36737 29600
rect 36771 29597 36783 29631
rect 36725 29591 36783 29597
rect 29086 29560 29092 29572
rect 25608 29532 29092 29560
rect 25510 29523 25568 29529
rect 29086 29520 29092 29532
rect 29144 29520 29150 29572
rect 31766 29563 31824 29569
rect 31766 29529 31778 29563
rect 31812 29529 31824 29563
rect 31766 29523 31824 29529
rect 35152 29563 35210 29569
rect 35152 29529 35164 29563
rect 35198 29560 35210 29563
rect 35434 29560 35440 29572
rect 35198 29532 35440 29560
rect 35198 29529 35210 29532
rect 35152 29523 35210 29529
rect 12621 29495 12679 29501
rect 12621 29461 12633 29495
rect 12667 29492 12679 29495
rect 12894 29492 12900 29504
rect 12667 29464 12900 29492
rect 12667 29461 12679 29464
rect 12621 29455 12679 29461
rect 12894 29452 12900 29464
rect 12952 29492 12958 29504
rect 13538 29492 13544 29504
rect 12952 29464 13544 29492
rect 12952 29452 12958 29464
rect 13538 29452 13544 29464
rect 13596 29452 13602 29504
rect 14274 29492 14280 29504
rect 14235 29464 14280 29492
rect 14274 29452 14280 29464
rect 14332 29452 14338 29504
rect 15197 29495 15255 29501
rect 15197 29461 15209 29495
rect 15243 29492 15255 29495
rect 15378 29492 15384 29504
rect 15243 29464 15384 29492
rect 15243 29461 15255 29464
rect 15197 29455 15255 29461
rect 15378 29452 15384 29464
rect 15436 29452 15442 29504
rect 15657 29495 15715 29501
rect 15657 29461 15669 29495
rect 15703 29492 15715 29495
rect 15746 29492 15752 29504
rect 15703 29464 15752 29492
rect 15703 29461 15715 29464
rect 15657 29455 15715 29461
rect 15746 29452 15752 29464
rect 15804 29452 15810 29504
rect 17218 29492 17224 29504
rect 17179 29464 17224 29492
rect 17218 29452 17224 29464
rect 17276 29452 17282 29504
rect 21177 29495 21235 29501
rect 21177 29461 21189 29495
rect 21223 29492 21235 29495
rect 22094 29492 22100 29504
rect 21223 29464 22100 29492
rect 21223 29461 21235 29464
rect 21177 29455 21235 29461
rect 22094 29452 22100 29464
rect 22152 29452 22158 29504
rect 22738 29492 22744 29504
rect 22699 29464 22744 29492
rect 22738 29452 22744 29464
rect 22796 29452 22802 29504
rect 24394 29492 24400 29504
rect 24355 29464 24400 29492
rect 24394 29452 24400 29464
rect 24452 29452 24458 29504
rect 28166 29452 28172 29504
rect 28224 29492 28230 29504
rect 30653 29495 30711 29501
rect 30653 29492 30665 29495
rect 28224 29464 30665 29492
rect 28224 29452 28230 29464
rect 30653 29461 30665 29464
rect 30699 29461 30711 29495
rect 31772 29492 31800 29523
rect 35434 29520 35440 29532
rect 35492 29520 35498 29572
rect 36538 29520 36544 29572
rect 36596 29560 36602 29572
rect 36970 29563 37028 29569
rect 36970 29560 36982 29563
rect 36596 29532 36982 29560
rect 36596 29520 36602 29532
rect 36970 29529 36982 29532
rect 37016 29529 37028 29563
rect 36970 29523 37028 29529
rect 31846 29492 31852 29504
rect 31772 29464 31852 29492
rect 30653 29455 30711 29461
rect 31846 29452 31852 29464
rect 31904 29452 31910 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 10134 29248 10140 29300
rect 10192 29288 10198 29300
rect 10229 29291 10287 29297
rect 10229 29288 10241 29291
rect 10192 29260 10241 29288
rect 10192 29248 10198 29260
rect 10229 29257 10241 29260
rect 10275 29257 10287 29291
rect 13170 29288 13176 29300
rect 13131 29260 13176 29288
rect 10229 29251 10287 29257
rect 13170 29248 13176 29260
rect 13228 29248 13234 29300
rect 15565 29291 15623 29297
rect 15565 29257 15577 29291
rect 15611 29288 15623 29291
rect 16298 29288 16304 29300
rect 15611 29260 16304 29288
rect 15611 29257 15623 29260
rect 15565 29251 15623 29257
rect 16298 29248 16304 29260
rect 16356 29248 16362 29300
rect 17218 29248 17224 29300
rect 17276 29288 17282 29300
rect 25590 29288 25596 29300
rect 17276 29260 22232 29288
rect 17276 29248 17282 29260
rect 20806 29220 20812 29232
rect 20767 29192 20812 29220
rect 20806 29180 20812 29192
rect 20864 29180 20870 29232
rect 20901 29223 20959 29229
rect 20901 29189 20913 29223
rect 20947 29220 20959 29223
rect 20990 29220 20996 29232
rect 20947 29192 20996 29220
rect 20947 29189 20959 29192
rect 20901 29183 20959 29189
rect 20990 29180 20996 29192
rect 21048 29180 21054 29232
rect 22204 29220 22232 29260
rect 22572 29260 25596 29288
rect 22572 29220 22600 29260
rect 25590 29248 25596 29260
rect 25648 29248 25654 29300
rect 22204 29192 22600 29220
rect 22738 29180 22744 29232
rect 22796 29220 22802 29232
rect 25510 29223 25568 29229
rect 25510 29220 25522 29223
rect 22796 29192 25522 29220
rect 22796 29180 22802 29192
rect 25510 29189 25522 29192
rect 25556 29189 25568 29223
rect 25510 29183 25568 29189
rect 32306 29180 32312 29232
rect 32364 29220 32370 29232
rect 32364 29192 34284 29220
rect 32364 29180 32370 29192
rect 12158 29152 12164 29164
rect 12119 29124 12164 29152
rect 12158 29112 12164 29124
rect 12216 29112 12222 29164
rect 12986 29152 12992 29164
rect 12947 29124 12992 29152
rect 12986 29112 12992 29124
rect 13044 29112 13050 29164
rect 15378 29152 15384 29164
rect 15339 29124 15384 29152
rect 15378 29112 15384 29124
rect 15436 29112 15442 29164
rect 19334 29112 19340 29164
rect 19392 29152 19398 29164
rect 19521 29155 19579 29161
rect 19521 29152 19533 29155
rect 19392 29124 19533 29152
rect 19392 29112 19398 29124
rect 19521 29121 19533 29124
rect 19567 29121 19579 29155
rect 21818 29152 21824 29164
rect 21779 29124 21824 29152
rect 19521 29115 19579 29121
rect 21818 29112 21824 29124
rect 21876 29112 21882 29164
rect 22002 29152 22008 29164
rect 21963 29124 22008 29152
rect 22002 29112 22008 29124
rect 22060 29112 22066 29164
rect 22189 29155 22247 29161
rect 22189 29121 22201 29155
rect 22235 29152 22247 29155
rect 22462 29152 22468 29164
rect 22235 29124 22468 29152
rect 22235 29121 22247 29124
rect 22189 29115 22247 29121
rect 22462 29112 22468 29124
rect 22520 29112 22526 29164
rect 29098 29155 29156 29161
rect 29098 29152 29110 29155
rect 24320 29124 29110 29152
rect 8570 29044 8576 29096
rect 8628 29084 8634 29096
rect 12526 29084 12532 29096
rect 8628 29056 12532 29084
rect 8628 29044 8634 29056
rect 12526 29044 12532 29056
rect 12584 29084 12590 29096
rect 13722 29084 13728 29096
rect 12584 29056 13728 29084
rect 12584 29044 12590 29056
rect 13722 29044 13728 29056
rect 13780 29044 13786 29096
rect 15194 29084 15200 29096
rect 15155 29056 15200 29084
rect 15194 29044 15200 29056
rect 15252 29044 15258 29096
rect 20717 29087 20775 29093
rect 20717 29053 20729 29087
rect 20763 29084 20775 29087
rect 21082 29084 21088 29096
rect 20763 29056 21088 29084
rect 20763 29053 20775 29056
rect 20717 29047 20775 29053
rect 21082 29044 21088 29056
rect 21140 29044 21146 29096
rect 21836 29084 21864 29112
rect 22649 29087 22707 29093
rect 22649 29084 22661 29087
rect 21836 29056 22661 29084
rect 22649 29053 22661 29056
rect 22695 29053 22707 29087
rect 22649 29047 22707 29053
rect 10502 28976 10508 29028
rect 10560 29016 10566 29028
rect 10781 29019 10839 29025
rect 10781 29016 10793 29019
rect 10560 28988 10793 29016
rect 10560 28976 10566 28988
rect 10781 28985 10793 28988
rect 10827 28985 10839 29019
rect 12342 29016 12348 29028
rect 12303 28988 12348 29016
rect 10781 28979 10839 28985
rect 12342 28976 12348 28988
rect 12400 28976 12406 29028
rect 15746 28976 15752 29028
rect 15804 29016 15810 29028
rect 16025 29019 16083 29025
rect 16025 29016 16037 29019
rect 15804 28988 16037 29016
rect 15804 28976 15810 28988
rect 16025 28985 16037 28988
rect 16071 28985 16083 29019
rect 16025 28979 16083 28985
rect 19705 29019 19763 29025
rect 19705 28985 19717 29019
rect 19751 29016 19763 29019
rect 24320 29016 24348 29124
rect 29098 29121 29110 29124
rect 29144 29121 29156 29155
rect 29098 29115 29156 29121
rect 29270 29112 29276 29164
rect 29328 29152 29334 29164
rect 29365 29155 29423 29161
rect 29365 29152 29377 29155
rect 29328 29124 29377 29152
rect 29328 29112 29334 29124
rect 29365 29121 29377 29124
rect 29411 29121 29423 29155
rect 29365 29115 29423 29121
rect 30558 29112 30564 29164
rect 30616 29152 30622 29164
rect 34256 29161 34284 29192
rect 33974 29155 34032 29161
rect 33974 29152 33986 29155
rect 30616 29124 33986 29152
rect 30616 29112 30622 29124
rect 33974 29121 33986 29124
rect 34020 29121 34032 29155
rect 33974 29115 34032 29121
rect 34241 29155 34299 29161
rect 34241 29121 34253 29155
rect 34287 29121 34299 29155
rect 34241 29115 34299 29121
rect 25777 29087 25835 29093
rect 25777 29053 25789 29087
rect 25823 29084 25835 29087
rect 26510 29084 26516 29096
rect 25823 29056 26516 29084
rect 25823 29053 25835 29056
rect 25777 29047 25835 29053
rect 26510 29044 26516 29056
rect 26568 29044 26574 29096
rect 19751 28988 24348 29016
rect 24397 29019 24455 29025
rect 19751 28985 19763 28988
rect 19705 28979 19763 28985
rect 24397 28985 24409 29019
rect 24443 29016 24455 29019
rect 24486 29016 24492 29028
rect 24443 28988 24492 29016
rect 24443 28985 24455 28988
rect 24397 28979 24455 28985
rect 24486 28976 24492 28988
rect 24544 28976 24550 29028
rect 27982 29016 27988 29028
rect 27943 28988 27988 29016
rect 27982 28976 27988 28988
rect 28040 28976 28046 29028
rect 32858 29016 32864 29028
rect 32819 28988 32864 29016
rect 32858 28976 32864 28988
rect 32916 28976 32922 29028
rect 9582 28908 9588 28960
rect 9640 28948 9646 28960
rect 9677 28951 9735 28957
rect 9677 28948 9689 28951
rect 9640 28920 9689 28948
rect 9640 28908 9646 28920
rect 9677 28917 9689 28920
rect 9723 28917 9735 28951
rect 9677 28911 9735 28917
rect 10870 28908 10876 28960
rect 10928 28948 10934 28960
rect 11517 28951 11575 28957
rect 11517 28948 11529 28951
rect 10928 28920 11529 28948
rect 10928 28908 10934 28920
rect 11517 28917 11529 28920
rect 11563 28917 11575 28951
rect 11517 28911 11575 28917
rect 21174 28908 21180 28960
rect 21232 28948 21238 28960
rect 21269 28951 21327 28957
rect 21269 28948 21281 28951
rect 21232 28920 21281 28948
rect 21232 28908 21238 28920
rect 21269 28917 21281 28920
rect 21315 28917 21327 28951
rect 21269 28911 21327 28917
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 14090 28744 14096 28756
rect 14051 28716 14096 28744
rect 14090 28704 14096 28716
rect 14148 28704 14154 28756
rect 17405 28747 17463 28753
rect 17405 28713 17417 28747
rect 17451 28744 17463 28747
rect 17494 28744 17500 28756
rect 17451 28716 17500 28744
rect 17451 28713 17463 28716
rect 17405 28707 17463 28713
rect 17494 28704 17500 28716
rect 17552 28704 17558 28756
rect 21818 28704 21824 28756
rect 21876 28744 21882 28756
rect 27617 28747 27675 28753
rect 27617 28744 27629 28747
rect 21876 28716 27629 28744
rect 21876 28704 21882 28716
rect 27617 28713 27629 28716
rect 27663 28713 27675 28747
rect 30929 28747 30987 28753
rect 30929 28744 30941 28747
rect 27617 28707 27675 28713
rect 27724 28716 30941 28744
rect 12066 28636 12072 28688
rect 12124 28676 12130 28688
rect 15654 28676 15660 28688
rect 12124 28648 15660 28676
rect 12124 28636 12130 28648
rect 15654 28636 15660 28648
rect 15712 28636 15718 28688
rect 18598 28636 18604 28688
rect 18656 28676 18662 28688
rect 25041 28679 25099 28685
rect 25041 28676 25053 28679
rect 18656 28648 25053 28676
rect 18656 28636 18662 28648
rect 25041 28645 25053 28648
rect 25087 28645 25099 28679
rect 25041 28639 25099 28645
rect 9582 28568 9588 28620
rect 9640 28608 9646 28620
rect 9677 28611 9735 28617
rect 9677 28608 9689 28611
rect 9640 28580 9689 28608
rect 9640 28568 9646 28580
rect 9677 28577 9689 28580
rect 9723 28608 9735 28611
rect 10781 28611 10839 28617
rect 10781 28608 10793 28611
rect 9723 28580 10793 28608
rect 9723 28577 9735 28580
rect 9677 28571 9735 28577
rect 10781 28577 10793 28580
rect 10827 28608 10839 28611
rect 15749 28611 15807 28617
rect 10827 28580 12940 28608
rect 10827 28577 10839 28580
rect 10781 28571 10839 28577
rect 5810 28500 5816 28552
rect 5868 28540 5874 28552
rect 5868 28512 6914 28540
rect 5868 28500 5874 28512
rect 6886 28472 6914 28512
rect 9122 28500 9128 28552
rect 9180 28540 9186 28552
rect 9493 28543 9551 28549
rect 9493 28540 9505 28543
rect 9180 28512 9505 28540
rect 9180 28500 9186 28512
rect 9493 28509 9505 28512
rect 9539 28540 9551 28543
rect 10502 28540 10508 28552
rect 9539 28512 10508 28540
rect 9539 28509 9551 28512
rect 9493 28503 9551 28509
rect 10502 28500 10508 28512
rect 10560 28500 10566 28552
rect 10689 28543 10747 28549
rect 10689 28509 10701 28543
rect 10735 28540 10747 28543
rect 10870 28540 10876 28552
rect 10735 28512 10876 28540
rect 10735 28509 10747 28512
rect 10689 28503 10747 28509
rect 10870 28500 10876 28512
rect 10928 28500 10934 28552
rect 11606 28540 11612 28552
rect 11567 28512 11612 28540
rect 11606 28500 11612 28512
rect 11664 28500 11670 28552
rect 10597 28475 10655 28481
rect 10597 28472 10609 28475
rect 6886 28444 10609 28472
rect 10597 28441 10609 28444
rect 10643 28472 10655 28475
rect 12342 28472 12348 28484
rect 10643 28444 12348 28472
rect 10643 28441 10655 28444
rect 10597 28435 10655 28441
rect 12342 28432 12348 28444
rect 12400 28432 12406 28484
rect 9030 28404 9036 28416
rect 8991 28376 9036 28404
rect 9030 28364 9036 28376
rect 9088 28364 9094 28416
rect 9401 28407 9459 28413
rect 9401 28373 9413 28407
rect 9447 28404 9459 28407
rect 10042 28404 10048 28416
rect 9447 28376 10048 28404
rect 9447 28373 9459 28376
rect 9401 28367 9459 28373
rect 10042 28364 10048 28376
rect 10100 28364 10106 28416
rect 10226 28404 10232 28416
rect 10187 28376 10232 28404
rect 10226 28364 10232 28376
rect 10284 28364 10290 28416
rect 11790 28404 11796 28416
rect 11751 28376 11796 28404
rect 11790 28364 11796 28376
rect 11848 28364 11854 28416
rect 12912 28413 12940 28580
rect 15749 28577 15761 28611
rect 15795 28608 15807 28611
rect 20530 28608 20536 28620
rect 15795 28580 20536 28608
rect 15795 28577 15807 28580
rect 15749 28571 15807 28577
rect 14274 28540 14280 28552
rect 14235 28512 14280 28540
rect 14274 28500 14280 28512
rect 14332 28500 14338 28552
rect 14461 28543 14519 28549
rect 14461 28509 14473 28543
rect 14507 28540 14519 28543
rect 14507 28512 15240 28540
rect 14507 28509 14519 28512
rect 14461 28503 14519 28509
rect 15212 28484 15240 28512
rect 15010 28472 15016 28484
rect 14923 28444 15016 28472
rect 15010 28432 15016 28444
rect 15068 28432 15074 28484
rect 15194 28472 15200 28484
rect 15155 28444 15200 28472
rect 15194 28432 15200 28444
rect 15252 28432 15258 28484
rect 12897 28407 12955 28413
rect 12897 28373 12909 28407
rect 12943 28404 12955 28407
rect 13814 28404 13820 28416
rect 12943 28376 13820 28404
rect 12943 28373 12955 28376
rect 12897 28367 12955 28373
rect 13814 28364 13820 28376
rect 13872 28364 13878 28416
rect 15028 28404 15056 28432
rect 15764 28404 15792 28571
rect 20530 28568 20536 28580
rect 20588 28568 20594 28620
rect 21082 28568 21088 28620
rect 21140 28608 21146 28620
rect 21818 28608 21824 28620
rect 21140 28580 21824 28608
rect 21140 28568 21146 28580
rect 21818 28568 21824 28580
rect 21876 28568 21882 28620
rect 27724 28608 27752 28716
rect 30929 28713 30941 28716
rect 30975 28713 30987 28747
rect 30929 28707 30987 28713
rect 38010 28704 38016 28756
rect 38068 28744 38074 28756
rect 38105 28747 38163 28753
rect 38105 28744 38117 28747
rect 38068 28716 38117 28744
rect 38068 28704 38074 28716
rect 38105 28713 38117 28716
rect 38151 28713 38163 28747
rect 38105 28707 38163 28713
rect 26344 28580 27752 28608
rect 28997 28611 29055 28617
rect 17037 28543 17095 28549
rect 17037 28509 17049 28543
rect 17083 28509 17095 28543
rect 17218 28540 17224 28552
rect 17179 28512 17224 28540
rect 17037 28503 17095 28509
rect 17052 28472 17080 28503
rect 17218 28500 17224 28512
rect 17276 28500 17282 28552
rect 21174 28540 21180 28552
rect 21135 28512 21180 28540
rect 21174 28500 21180 28512
rect 21232 28500 21238 28552
rect 26344 28540 26372 28580
rect 28997 28577 29009 28611
rect 29043 28608 29055 28611
rect 29270 28608 29276 28620
rect 29043 28580 29276 28608
rect 29043 28577 29055 28580
rect 28997 28571 29055 28577
rect 29270 28568 29276 28580
rect 29328 28568 29334 28620
rect 32306 28608 32312 28620
rect 32267 28580 32312 28608
rect 32306 28568 32312 28580
rect 32364 28568 32370 28620
rect 21284 28512 26372 28540
rect 26421 28543 26479 28549
rect 18782 28472 18788 28484
rect 17052 28444 18788 28472
rect 18782 28432 18788 28444
rect 18840 28432 18846 28484
rect 18874 28432 18880 28484
rect 18932 28472 18938 28484
rect 21284 28472 21312 28512
rect 26421 28509 26433 28543
rect 26467 28540 26479 28543
rect 26510 28540 26516 28552
rect 26467 28512 26516 28540
rect 26467 28509 26479 28512
rect 26421 28503 26479 28509
rect 26510 28500 26516 28512
rect 26568 28500 26574 28552
rect 36725 28543 36783 28549
rect 36725 28509 36737 28543
rect 36771 28540 36783 28543
rect 36814 28540 36820 28552
rect 36771 28512 36820 28540
rect 36771 28509 36783 28512
rect 36725 28503 36783 28509
rect 36814 28500 36820 28512
rect 36872 28500 36878 28552
rect 18932 28444 21312 28472
rect 21376 28444 25452 28472
rect 18932 28432 18938 28444
rect 16206 28404 16212 28416
rect 15028 28376 15792 28404
rect 16167 28376 16212 28404
rect 16206 28364 16212 28376
rect 16264 28364 16270 28416
rect 21376 28413 21404 28444
rect 21361 28407 21419 28413
rect 21361 28373 21373 28407
rect 21407 28373 21419 28407
rect 25424 28404 25452 28444
rect 25590 28432 25596 28484
rect 25648 28472 25654 28484
rect 26154 28475 26212 28481
rect 26154 28472 26166 28475
rect 25648 28444 26166 28472
rect 25648 28432 25654 28444
rect 26154 28441 26166 28444
rect 26200 28441 26212 28475
rect 28730 28475 28788 28481
rect 28730 28472 28742 28475
rect 26154 28435 26212 28441
rect 26252 28444 28742 28472
rect 26252 28404 26280 28444
rect 28730 28441 28742 28444
rect 28776 28441 28788 28475
rect 28730 28435 28788 28441
rect 31754 28432 31760 28484
rect 31812 28472 31818 28484
rect 32042 28475 32100 28481
rect 32042 28472 32054 28475
rect 31812 28444 32054 28472
rect 31812 28432 31818 28444
rect 32042 28441 32054 28444
rect 32088 28441 32100 28475
rect 32042 28435 32100 28441
rect 36170 28432 36176 28484
rect 36228 28472 36234 28484
rect 36970 28475 37028 28481
rect 36970 28472 36982 28475
rect 36228 28444 36982 28472
rect 36228 28432 36234 28444
rect 36970 28441 36982 28444
rect 37016 28441 37028 28475
rect 36970 28435 37028 28441
rect 25424 28376 26280 28404
rect 21361 28367 21419 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 9950 28200 9956 28212
rect 9911 28172 9956 28200
rect 9950 28160 9956 28172
rect 10008 28160 10014 28212
rect 12158 28160 12164 28212
rect 12216 28200 12222 28212
rect 12253 28203 12311 28209
rect 12253 28200 12265 28203
rect 12216 28172 12265 28200
rect 12216 28160 12222 28172
rect 12253 28169 12265 28172
rect 12299 28169 12311 28203
rect 12253 28163 12311 28169
rect 12713 28203 12771 28209
rect 12713 28169 12725 28203
rect 12759 28200 12771 28203
rect 12986 28200 12992 28212
rect 12759 28172 12992 28200
rect 12759 28169 12771 28172
rect 12713 28163 12771 28169
rect 12986 28160 12992 28172
rect 13044 28160 13050 28212
rect 15286 28160 15292 28212
rect 15344 28200 15350 28212
rect 15381 28203 15439 28209
rect 15381 28200 15393 28203
rect 15344 28172 15393 28200
rect 15344 28160 15350 28172
rect 15381 28169 15393 28172
rect 15427 28169 15439 28203
rect 15381 28163 15439 28169
rect 15654 28160 15660 28212
rect 15712 28200 15718 28212
rect 15749 28203 15807 28209
rect 15749 28200 15761 28203
rect 15712 28172 15761 28200
rect 15712 28160 15718 28172
rect 15749 28169 15761 28172
rect 15795 28169 15807 28203
rect 15749 28163 15807 28169
rect 19153 28203 19211 28209
rect 19153 28169 19165 28203
rect 19199 28200 19211 28203
rect 19334 28200 19340 28212
rect 19199 28172 19340 28200
rect 19199 28169 19211 28172
rect 19153 28163 19211 28169
rect 19334 28160 19340 28172
rect 19392 28160 19398 28212
rect 11790 28092 11796 28144
rect 11848 28132 11854 28144
rect 25142 28135 25200 28141
rect 25142 28132 25154 28135
rect 11848 28104 25154 28132
rect 11848 28092 11854 28104
rect 25142 28101 25154 28104
rect 25188 28101 25200 28135
rect 25142 28095 25200 28101
rect 29270 28092 29276 28144
rect 29328 28132 29334 28144
rect 29328 28104 30052 28132
rect 29328 28092 29334 28104
rect 9030 28064 9036 28076
rect 8991 28036 9036 28064
rect 9030 28024 9036 28036
rect 9088 28024 9094 28076
rect 9217 28067 9275 28073
rect 9217 28033 9229 28067
rect 9263 28064 9275 28067
rect 9769 28067 9827 28073
rect 9769 28064 9781 28067
rect 9263 28036 9781 28064
rect 9263 28033 9275 28036
rect 9217 28027 9275 28033
rect 9769 28033 9781 28036
rect 9815 28033 9827 28067
rect 9769 28027 9827 28033
rect 10226 28024 10232 28076
rect 10284 28064 10290 28076
rect 10597 28067 10655 28073
rect 10597 28064 10609 28067
rect 10284 28036 10609 28064
rect 10284 28024 10290 28036
rect 10597 28033 10609 28036
rect 10643 28033 10655 28067
rect 11882 28064 11888 28076
rect 11843 28036 11888 28064
rect 10597 28027 10655 28033
rect 11882 28024 11888 28036
rect 11940 28024 11946 28076
rect 12066 28064 12072 28076
rect 12027 28036 12072 28064
rect 12066 28024 12072 28036
rect 12124 28024 12130 28076
rect 12897 28067 12955 28073
rect 12897 28033 12909 28067
rect 12943 28064 12955 28067
rect 13262 28064 13268 28076
rect 12943 28036 13268 28064
rect 12943 28033 12955 28036
rect 12897 28027 12955 28033
rect 13262 28024 13268 28036
rect 13320 28024 13326 28076
rect 15841 28067 15899 28073
rect 15841 28033 15853 28067
rect 15887 28064 15899 28067
rect 16206 28064 16212 28076
rect 15887 28036 16212 28064
rect 15887 28033 15899 28036
rect 15841 28027 15899 28033
rect 16206 28024 16212 28036
rect 16264 28024 16270 28076
rect 16666 28064 16672 28076
rect 16627 28036 16672 28064
rect 16666 28024 16672 28036
rect 16724 28024 16730 28076
rect 18966 28064 18972 28076
rect 18927 28036 18972 28064
rect 18966 28024 18972 28036
rect 19024 28024 19030 28076
rect 29730 28064 29736 28076
rect 29788 28073 29794 28076
rect 30024 28073 30052 28104
rect 34514 28092 34520 28144
rect 34572 28132 34578 28144
rect 35170 28135 35228 28141
rect 35170 28132 35182 28135
rect 34572 28104 35182 28132
rect 34572 28092 34578 28104
rect 35170 28101 35182 28104
rect 35216 28101 35228 28135
rect 35170 28095 35228 28101
rect 29700 28036 29736 28064
rect 29730 28024 29736 28036
rect 29788 28027 29800 28073
rect 30009 28067 30067 28073
rect 30009 28033 30021 28067
rect 30055 28033 30067 28067
rect 30009 28027 30067 28033
rect 29788 28024 29794 28027
rect 8849 27999 8907 28005
rect 8849 27965 8861 27999
rect 8895 27996 8907 27999
rect 10413 27999 10471 28005
rect 10413 27996 10425 27999
rect 8895 27968 10425 27996
rect 8895 27965 8907 27968
rect 8849 27959 8907 27965
rect 10413 27965 10425 27968
rect 10459 27996 10471 27999
rect 11054 27996 11060 28008
rect 10459 27968 11060 27996
rect 10459 27965 10471 27968
rect 10413 27959 10471 27965
rect 11054 27956 11060 27968
rect 11112 27996 11118 28008
rect 11900 27996 11928 28024
rect 11112 27968 11928 27996
rect 13081 27999 13139 28005
rect 11112 27956 11118 27968
rect 13081 27965 13093 27999
rect 13127 27996 13139 27999
rect 15194 27996 15200 28008
rect 13127 27968 15200 27996
rect 13127 27965 13139 27968
rect 13081 27959 13139 27965
rect 15194 27956 15200 27968
rect 15252 27956 15258 28008
rect 15930 27996 15936 28008
rect 15891 27968 15936 27996
rect 15930 27956 15936 27968
rect 15988 27956 15994 28008
rect 18782 27996 18788 28008
rect 18743 27968 18788 27996
rect 18782 27956 18788 27968
rect 18840 27956 18846 28008
rect 25409 27999 25467 28005
rect 25409 27965 25421 27999
rect 25455 27996 25467 27999
rect 26234 27996 26240 28008
rect 25455 27968 26240 27996
rect 25455 27965 25467 27968
rect 25409 27959 25467 27965
rect 26234 27956 26240 27968
rect 26292 27996 26298 28008
rect 26510 27996 26516 28008
rect 26292 27968 26516 27996
rect 26292 27956 26298 27968
rect 26510 27956 26516 27968
rect 26568 27956 26574 28008
rect 35437 27999 35495 28005
rect 35437 27965 35449 27999
rect 35483 27996 35495 27999
rect 35894 27996 35900 28008
rect 35483 27968 35900 27996
rect 35483 27965 35495 27968
rect 35437 27959 35495 27965
rect 35894 27956 35900 27968
rect 35952 27996 35958 28008
rect 36998 27996 37004 28008
rect 35952 27968 37004 27996
rect 35952 27956 35958 27968
rect 36998 27956 37004 27968
rect 37056 27956 37062 28008
rect 13446 27888 13452 27940
rect 13504 27928 13510 27940
rect 16850 27928 16856 27940
rect 13504 27900 15056 27928
rect 16811 27900 16856 27928
rect 13504 27888 13510 27900
rect 10781 27863 10839 27869
rect 10781 27829 10793 27863
rect 10827 27860 10839 27863
rect 11698 27860 11704 27872
rect 10827 27832 11704 27860
rect 10827 27829 10839 27832
rect 10781 27823 10839 27829
rect 11698 27820 11704 27832
rect 11756 27820 11762 27872
rect 13538 27860 13544 27872
rect 13499 27832 13544 27860
rect 13538 27820 13544 27832
rect 13596 27820 13602 27872
rect 14918 27860 14924 27872
rect 14879 27832 14924 27860
rect 14918 27820 14924 27832
rect 14976 27820 14982 27872
rect 15028 27860 15056 27900
rect 16850 27888 16856 27900
rect 16908 27888 16914 27940
rect 24029 27931 24087 27937
rect 24029 27928 24041 27931
rect 16960 27900 24041 27928
rect 16960 27860 16988 27900
rect 24029 27897 24041 27900
rect 24075 27897 24087 27931
rect 24029 27891 24087 27897
rect 15028 27832 16988 27860
rect 20257 27863 20315 27869
rect 20257 27829 20269 27863
rect 20303 27860 20315 27863
rect 20530 27860 20536 27872
rect 20303 27832 20536 27860
rect 20303 27829 20315 27832
rect 20257 27823 20315 27829
rect 20530 27820 20536 27832
rect 20588 27820 20594 27872
rect 25038 27820 25044 27872
rect 25096 27860 25102 27872
rect 28629 27863 28687 27869
rect 28629 27860 28641 27863
rect 25096 27832 28641 27860
rect 25096 27820 25102 27832
rect 28629 27829 28641 27832
rect 28675 27829 28687 27863
rect 28629 27823 28687 27829
rect 32030 27820 32036 27872
rect 32088 27860 32094 27872
rect 34057 27863 34115 27869
rect 34057 27860 34069 27863
rect 32088 27832 34069 27860
rect 32088 27820 32094 27832
rect 34057 27829 34069 27832
rect 34103 27829 34115 27863
rect 34057 27823 34115 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 11054 27656 11060 27668
rect 10888 27628 11060 27656
rect 10888 27529 10916 27628
rect 11054 27616 11060 27628
rect 11112 27616 11118 27668
rect 11241 27659 11299 27665
rect 11241 27625 11253 27659
rect 11287 27656 11299 27659
rect 11606 27656 11612 27668
rect 11287 27628 11612 27656
rect 11287 27625 11299 27628
rect 11241 27619 11299 27625
rect 11606 27616 11612 27628
rect 11664 27616 11670 27668
rect 11977 27659 12035 27665
rect 11977 27625 11989 27659
rect 12023 27656 12035 27659
rect 12066 27656 12072 27668
rect 12023 27628 12072 27656
rect 12023 27625 12035 27628
rect 11977 27619 12035 27625
rect 12066 27616 12072 27628
rect 12124 27616 12130 27668
rect 24872 27628 25820 27656
rect 15657 27591 15715 27597
rect 15657 27557 15669 27591
rect 15703 27588 15715 27591
rect 16666 27588 16672 27600
rect 15703 27560 16672 27588
rect 15703 27557 15715 27560
rect 15657 27551 15715 27557
rect 16666 27548 16672 27560
rect 16724 27548 16730 27600
rect 18049 27591 18107 27597
rect 18049 27557 18061 27591
rect 18095 27557 18107 27591
rect 18690 27588 18696 27600
rect 18651 27560 18696 27588
rect 18049 27551 18107 27557
rect 10873 27523 10931 27529
rect 10873 27489 10885 27523
rect 10919 27489 10931 27523
rect 10873 27483 10931 27489
rect 12621 27523 12679 27529
rect 12621 27489 12633 27523
rect 12667 27520 12679 27523
rect 12802 27520 12808 27532
rect 12667 27492 12808 27520
rect 12667 27489 12679 27492
rect 12621 27483 12679 27489
rect 12802 27480 12808 27492
rect 12860 27480 12866 27532
rect 13814 27480 13820 27532
rect 13872 27520 13878 27532
rect 14277 27523 14335 27529
rect 14277 27520 14289 27523
rect 13872 27492 14289 27520
rect 13872 27480 13878 27492
rect 14277 27489 14289 27492
rect 14323 27520 14335 27523
rect 14918 27520 14924 27532
rect 14323 27492 14924 27520
rect 14323 27489 14335 27492
rect 14277 27483 14335 27489
rect 14918 27480 14924 27492
rect 14976 27480 14982 27532
rect 15194 27480 15200 27532
rect 15252 27520 15258 27532
rect 15289 27523 15347 27529
rect 15289 27520 15301 27523
rect 15252 27492 15301 27520
rect 15252 27480 15258 27492
rect 15289 27489 15301 27492
rect 15335 27520 15347 27523
rect 16482 27520 16488 27532
rect 15335 27492 16488 27520
rect 15335 27489 15347 27492
rect 15289 27483 15347 27489
rect 16482 27480 16488 27492
rect 16540 27480 16546 27532
rect 18064 27520 18092 27551
rect 18690 27548 18696 27560
rect 18748 27548 18754 27600
rect 19242 27588 19248 27600
rect 19203 27560 19248 27588
rect 19242 27548 19248 27560
rect 19300 27548 19306 27600
rect 24872 27588 24900 27628
rect 20088 27560 24900 27588
rect 25792 27588 25820 27628
rect 33244 27628 34192 27656
rect 25792 27560 26556 27588
rect 20088 27520 20116 27560
rect 18064 27492 20116 27520
rect 20717 27523 20775 27529
rect 20717 27489 20729 27523
rect 20763 27520 20775 27523
rect 26418 27520 26424 27532
rect 20763 27492 22094 27520
rect 20763 27489 20775 27492
rect 20717 27483 20775 27489
rect 11054 27452 11060 27464
rect 11015 27424 11060 27452
rect 11054 27412 11060 27424
rect 11112 27412 11118 27464
rect 11146 27412 11152 27464
rect 11204 27452 11210 27464
rect 12345 27455 12403 27461
rect 12345 27452 12357 27455
rect 11204 27424 12357 27452
rect 11204 27412 11210 27424
rect 12345 27421 12357 27424
rect 12391 27452 12403 27455
rect 13265 27455 13323 27461
rect 13265 27452 13277 27455
rect 12391 27424 13277 27452
rect 12391 27421 12403 27424
rect 12345 27415 12403 27421
rect 13265 27421 13277 27424
rect 13311 27452 13323 27455
rect 15470 27452 15476 27464
rect 13311 27424 15332 27452
rect 15431 27424 15476 27452
rect 13311 27421 13323 27424
rect 13265 27415 13323 27421
rect 10502 27344 10508 27396
rect 10560 27384 10566 27396
rect 12437 27387 12495 27393
rect 12437 27384 12449 27387
rect 10560 27356 12449 27384
rect 10560 27344 10566 27356
rect 12437 27353 12449 27356
rect 12483 27384 12495 27387
rect 13538 27384 13544 27396
rect 12483 27356 13544 27384
rect 12483 27353 12495 27356
rect 12437 27347 12495 27353
rect 13538 27344 13544 27356
rect 13596 27344 13602 27396
rect 14369 27387 14427 27393
rect 14369 27353 14381 27387
rect 14415 27384 14427 27387
rect 15194 27384 15200 27396
rect 14415 27356 15200 27384
rect 14415 27353 14427 27356
rect 14369 27347 14427 27353
rect 15194 27344 15200 27356
rect 15252 27344 15258 27396
rect 7558 27276 7564 27328
rect 7616 27316 7622 27328
rect 14458 27316 14464 27328
rect 7616 27288 14464 27316
rect 7616 27276 7622 27288
rect 14458 27276 14464 27288
rect 14516 27276 14522 27328
rect 14550 27276 14556 27328
rect 14608 27316 14614 27328
rect 14829 27319 14887 27325
rect 14829 27316 14841 27319
rect 14608 27288 14841 27316
rect 14608 27276 14614 27288
rect 14829 27285 14841 27288
rect 14875 27285 14887 27319
rect 15304 27316 15332 27424
rect 15470 27412 15476 27424
rect 15528 27412 15534 27464
rect 15654 27412 15660 27464
rect 15712 27452 15718 27464
rect 16393 27455 16451 27461
rect 16393 27452 16405 27455
rect 15712 27424 16405 27452
rect 15712 27412 15718 27424
rect 16393 27421 16405 27424
rect 16439 27421 16451 27455
rect 16393 27415 16451 27421
rect 17126 27412 17132 27464
rect 17184 27452 17190 27464
rect 17865 27455 17923 27461
rect 17865 27452 17877 27455
rect 17184 27424 17877 27452
rect 17184 27412 17190 27424
rect 17865 27421 17877 27424
rect 17911 27421 17923 27455
rect 18506 27452 18512 27464
rect 18467 27424 18512 27452
rect 17865 27415 17923 27421
rect 18506 27412 18512 27424
rect 18564 27412 18570 27464
rect 20349 27455 20407 27461
rect 20349 27421 20361 27455
rect 20395 27421 20407 27455
rect 20349 27415 20407 27421
rect 20533 27455 20591 27461
rect 20533 27421 20545 27455
rect 20579 27421 20591 27455
rect 20533 27415 20591 27421
rect 17862 27316 17868 27328
rect 15304 27288 17868 27316
rect 14829 27279 14887 27285
rect 17862 27276 17868 27288
rect 17920 27276 17926 27328
rect 19889 27319 19947 27325
rect 19889 27285 19901 27319
rect 19935 27316 19947 27319
rect 20364 27316 20392 27415
rect 20548 27384 20576 27415
rect 20806 27412 20812 27464
rect 20864 27452 20870 27464
rect 21637 27455 21695 27461
rect 21637 27452 21649 27455
rect 20864 27424 21649 27452
rect 20864 27412 20870 27424
rect 21637 27421 21649 27424
rect 21683 27421 21695 27455
rect 22066 27452 22094 27492
rect 25700 27492 26424 27520
rect 22281 27455 22339 27461
rect 22281 27452 22293 27455
rect 22066 27424 22293 27452
rect 21637 27415 21695 27421
rect 22281 27421 22293 27424
rect 22327 27421 22339 27455
rect 22281 27415 22339 27421
rect 22554 27412 22560 27464
rect 22612 27452 22618 27464
rect 25700 27452 25728 27492
rect 26418 27480 26424 27492
rect 26476 27480 26482 27532
rect 22612 27424 25728 27452
rect 25777 27455 25835 27461
rect 22612 27412 22618 27424
rect 25777 27421 25789 27455
rect 25823 27452 25835 27455
rect 26234 27452 26240 27464
rect 25823 27424 26240 27452
rect 25823 27421 25835 27424
rect 25777 27415 25835 27421
rect 26234 27412 26240 27424
rect 26292 27412 26298 27464
rect 26528 27452 26556 27560
rect 30098 27548 30104 27600
rect 30156 27588 30162 27600
rect 32769 27591 32827 27597
rect 32769 27588 32781 27591
rect 30156 27560 32781 27588
rect 30156 27548 30162 27560
rect 32769 27557 32781 27560
rect 32815 27557 32827 27591
rect 33244 27588 33272 27628
rect 32769 27551 32827 27557
rect 32876 27560 33272 27588
rect 34164 27588 34192 27628
rect 35621 27591 35679 27597
rect 35621 27588 35633 27591
rect 34164 27560 35633 27588
rect 27709 27523 27767 27529
rect 27709 27489 27721 27523
rect 27755 27520 27767 27523
rect 29270 27520 29276 27532
rect 27755 27492 29276 27520
rect 27755 27489 27767 27492
rect 27709 27483 27767 27489
rect 29270 27480 29276 27492
rect 29328 27480 29334 27532
rect 29362 27480 29368 27532
rect 29420 27520 29426 27532
rect 30190 27520 30196 27532
rect 29420 27492 30196 27520
rect 29420 27480 29426 27492
rect 30190 27480 30196 27492
rect 30248 27520 30254 27532
rect 32876 27520 32904 27560
rect 35621 27557 35633 27560
rect 35667 27557 35679 27591
rect 35621 27551 35679 27557
rect 30248 27492 32904 27520
rect 30248 27480 30254 27492
rect 30650 27452 30656 27464
rect 26528 27424 30656 27452
rect 30650 27412 30656 27424
rect 30708 27412 30714 27464
rect 31754 27412 31760 27464
rect 31812 27452 31818 27464
rect 31938 27452 31944 27464
rect 31812 27424 31944 27452
rect 31812 27412 31818 27424
rect 31938 27412 31944 27424
rect 31996 27412 32002 27464
rect 32306 27412 32312 27464
rect 32364 27452 32370 27464
rect 33042 27452 33048 27464
rect 32364 27424 33048 27452
rect 32364 27412 32370 27424
rect 33042 27412 33048 27424
rect 33100 27452 33106 27464
rect 34149 27455 34207 27461
rect 34149 27452 34161 27455
rect 33100 27424 34161 27452
rect 33100 27412 33106 27424
rect 34149 27421 34161 27424
rect 34195 27421 34207 27455
rect 36998 27452 37004 27464
rect 36959 27424 37004 27452
rect 34149 27415 34207 27421
rect 36998 27412 37004 27424
rect 37056 27412 37062 27464
rect 20714 27384 20720 27396
rect 20548 27356 20720 27384
rect 20714 27344 20720 27356
rect 20772 27344 20778 27396
rect 24854 27344 24860 27396
rect 24912 27384 24918 27396
rect 25510 27387 25568 27393
rect 25510 27384 25522 27387
rect 24912 27356 25522 27384
rect 24912 27344 24918 27356
rect 25510 27353 25522 27356
rect 25556 27353 25568 27387
rect 25510 27347 25568 27353
rect 26418 27344 26424 27396
rect 26476 27384 26482 27396
rect 27442 27387 27500 27393
rect 27442 27384 27454 27387
rect 26476 27356 27454 27384
rect 26476 27344 26482 27356
rect 27442 27353 27454 27356
rect 27488 27353 27500 27387
rect 27442 27347 27500 27353
rect 30742 27344 30748 27396
rect 30800 27384 30806 27396
rect 33882 27387 33940 27393
rect 33882 27384 33894 27387
rect 30800 27356 33894 27384
rect 30800 27344 30806 27356
rect 33882 27353 33894 27356
rect 33928 27353 33940 27387
rect 36734 27387 36792 27393
rect 36734 27384 36746 27387
rect 33882 27347 33940 27353
rect 33980 27356 36746 27384
rect 20530 27316 20536 27328
rect 19935 27288 20536 27316
rect 19935 27285 19947 27288
rect 19889 27279 19947 27285
rect 20530 27276 20536 27288
rect 20588 27276 20594 27328
rect 21818 27316 21824 27328
rect 21779 27288 21824 27316
rect 21818 27276 21824 27288
rect 21876 27276 21882 27328
rect 22465 27319 22523 27325
rect 22465 27285 22477 27319
rect 22511 27316 22523 27319
rect 24302 27316 24308 27328
rect 22511 27288 24308 27316
rect 22511 27285 22523 27288
rect 22465 27279 22523 27285
rect 24302 27276 24308 27288
rect 24360 27276 24366 27328
rect 24394 27276 24400 27328
rect 24452 27316 24458 27328
rect 24452 27288 24497 27316
rect 24452 27276 24458 27288
rect 25038 27276 25044 27328
rect 25096 27316 25102 27328
rect 26329 27319 26387 27325
rect 26329 27316 26341 27319
rect 25096 27288 26341 27316
rect 25096 27276 25102 27288
rect 26329 27285 26341 27288
rect 26375 27285 26387 27319
rect 26329 27279 26387 27285
rect 30466 27276 30472 27328
rect 30524 27316 30530 27328
rect 33980 27316 34008 27356
rect 36734 27353 36746 27356
rect 36780 27353 36792 27387
rect 36734 27347 36792 27353
rect 30524 27288 34008 27316
rect 30524 27276 30530 27288
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 12250 27072 12256 27124
rect 12308 27112 12314 27124
rect 12345 27115 12403 27121
rect 12345 27112 12357 27115
rect 12308 27084 12357 27112
rect 12308 27072 12314 27084
rect 12345 27081 12357 27084
rect 12391 27081 12403 27115
rect 12345 27075 12403 27081
rect 12526 27072 12532 27124
rect 12584 27112 12590 27124
rect 12713 27115 12771 27121
rect 12713 27112 12725 27115
rect 12584 27084 12725 27112
rect 12584 27072 12590 27084
rect 12713 27081 12725 27084
rect 12759 27112 12771 27115
rect 13541 27115 13599 27121
rect 13541 27112 13553 27115
rect 12759 27084 13553 27112
rect 12759 27081 12771 27084
rect 12713 27075 12771 27081
rect 13541 27081 13553 27084
rect 13587 27081 13599 27115
rect 13541 27075 13599 27081
rect 17773 27115 17831 27121
rect 17773 27081 17785 27115
rect 17819 27112 17831 27115
rect 18506 27112 18512 27124
rect 17819 27084 18512 27112
rect 17819 27081 17831 27084
rect 17773 27075 17831 27081
rect 18506 27072 18512 27084
rect 18564 27072 18570 27124
rect 20806 27112 20812 27124
rect 20767 27084 20812 27112
rect 20806 27072 20812 27084
rect 20864 27072 20870 27124
rect 21818 27072 21824 27124
rect 21876 27112 21882 27124
rect 31478 27112 31484 27124
rect 21876 27084 31484 27112
rect 21876 27072 21882 27084
rect 31478 27072 31484 27084
rect 31536 27072 31542 27124
rect 32125 27115 32183 27121
rect 32125 27112 32137 27115
rect 31726 27084 32137 27112
rect 31726 27056 31754 27084
rect 32125 27081 32137 27084
rect 32171 27081 32183 27115
rect 35342 27112 35348 27124
rect 35303 27084 35348 27112
rect 32125 27075 32183 27081
rect 35342 27072 35348 27084
rect 35400 27112 35406 27124
rect 35618 27112 35624 27124
rect 35400 27084 35624 27112
rect 35400 27072 35406 27084
rect 35618 27072 35624 27084
rect 35676 27072 35682 27124
rect 14458 27004 14464 27056
rect 14516 27044 14522 27056
rect 15289 27047 15347 27053
rect 15289 27044 15301 27047
rect 14516 27016 15301 27044
rect 14516 27004 14522 27016
rect 15289 27013 15301 27016
rect 15335 27044 15347 27047
rect 15335 27016 17724 27044
rect 15335 27013 15347 27016
rect 15289 27007 15347 27013
rect 8570 26976 8576 26988
rect 8531 26948 8576 26976
rect 8570 26936 8576 26948
rect 8628 26936 8634 26988
rect 9122 26936 9128 26988
rect 9180 26976 9186 26988
rect 9401 26979 9459 26985
rect 9401 26976 9413 26979
rect 9180 26948 9413 26976
rect 9180 26936 9186 26948
rect 9401 26945 9413 26948
rect 9447 26945 9459 26979
rect 9401 26939 9459 26945
rect 9585 26979 9643 26985
rect 9585 26945 9597 26979
rect 9631 26976 9643 26979
rect 10045 26979 10103 26985
rect 10045 26976 10057 26979
rect 9631 26948 10057 26976
rect 9631 26945 9643 26948
rect 9585 26939 9643 26945
rect 10045 26945 10057 26948
rect 10091 26945 10103 26979
rect 10045 26939 10103 26945
rect 11238 26936 11244 26988
rect 11296 26976 11302 26988
rect 11609 26979 11667 26985
rect 11609 26976 11621 26979
rect 11296 26948 11621 26976
rect 11296 26936 11302 26948
rect 11609 26945 11621 26948
rect 11655 26945 11667 26979
rect 11609 26939 11667 26945
rect 12805 26979 12863 26985
rect 12805 26945 12817 26979
rect 12851 26976 12863 26979
rect 13170 26976 13176 26988
rect 12851 26948 13176 26976
rect 12851 26945 12863 26948
rect 12805 26939 12863 26945
rect 13170 26936 13176 26948
rect 13228 26936 13234 26988
rect 14366 26976 14372 26988
rect 14327 26948 14372 26976
rect 14366 26936 14372 26948
rect 14424 26936 14430 26988
rect 14550 26976 14556 26988
rect 14511 26948 14556 26976
rect 14550 26936 14556 26948
rect 14608 26936 14614 26988
rect 14918 26936 14924 26988
rect 14976 26976 14982 26988
rect 16942 26976 16948 26988
rect 14976 26948 16948 26976
rect 14976 26936 14982 26948
rect 16942 26936 16948 26948
rect 17000 26936 17006 26988
rect 17586 26976 17592 26988
rect 17547 26948 17592 26976
rect 17586 26936 17592 26948
rect 17644 26936 17650 26988
rect 17696 26976 17724 27016
rect 17862 27004 17868 27056
rect 17920 27044 17926 27056
rect 22554 27044 22560 27056
rect 17920 27016 22560 27044
rect 17920 27004 17926 27016
rect 22554 27004 22560 27016
rect 22612 27004 22618 27056
rect 22646 27004 22652 27056
rect 22704 27044 22710 27056
rect 29978 27047 30036 27053
rect 29978 27044 29990 27047
rect 22704 27016 29990 27044
rect 22704 27004 22710 27016
rect 29978 27013 29990 27016
rect 30024 27013 30036 27047
rect 29978 27007 30036 27013
rect 31110 27004 31116 27056
rect 31168 27044 31174 27056
rect 31662 27044 31668 27056
rect 31168 27016 31668 27044
rect 31168 27004 31174 27016
rect 31662 27004 31668 27016
rect 31720 27016 31754 27056
rect 31720 27004 31726 27016
rect 33042 27004 33048 27056
rect 33100 27044 33106 27056
rect 33100 27016 33548 27044
rect 33100 27004 33106 27016
rect 18138 26976 18144 26988
rect 17696 26948 18144 26976
rect 18138 26936 18144 26948
rect 18196 26936 18202 26988
rect 18782 26936 18788 26988
rect 18840 26976 18846 26988
rect 18877 26979 18935 26985
rect 18877 26976 18889 26979
rect 18840 26948 18889 26976
rect 18840 26936 18846 26948
rect 18877 26945 18889 26948
rect 18923 26945 18935 26979
rect 18877 26939 18935 26945
rect 19061 26979 19119 26985
rect 19061 26945 19073 26979
rect 19107 26945 19119 26979
rect 19061 26939 19119 26945
rect 19245 26979 19303 26985
rect 19245 26945 19257 26979
rect 19291 26976 19303 26979
rect 19705 26979 19763 26985
rect 19705 26976 19717 26979
rect 19291 26948 19717 26976
rect 19291 26945 19303 26948
rect 19245 26939 19303 26945
rect 19705 26945 19717 26948
rect 19751 26945 19763 26979
rect 20530 26976 20536 26988
rect 20491 26948 20536 26976
rect 19705 26939 19763 26945
rect 8389 26911 8447 26917
rect 8389 26877 8401 26911
rect 8435 26908 8447 26911
rect 9217 26911 9275 26917
rect 9217 26908 9229 26911
rect 8435 26880 9229 26908
rect 8435 26877 8447 26880
rect 8389 26871 8447 26877
rect 9217 26877 9229 26880
rect 9263 26908 9275 26911
rect 10962 26908 10968 26920
rect 9263 26880 10968 26908
rect 9263 26877 9275 26880
rect 9217 26871 9275 26877
rect 10962 26868 10968 26880
rect 11020 26868 11026 26920
rect 12894 26908 12900 26920
rect 12855 26880 12900 26908
rect 12894 26868 12900 26880
rect 12952 26868 12958 26920
rect 16482 26868 16488 26920
rect 16540 26908 16546 26920
rect 17405 26911 17463 26917
rect 17405 26908 17417 26911
rect 16540 26880 17417 26908
rect 16540 26868 16546 26880
rect 17405 26877 17417 26880
rect 17451 26908 17463 26911
rect 18800 26908 18828 26936
rect 17451 26880 18828 26908
rect 19076 26908 19104 26939
rect 20530 26936 20536 26948
rect 20588 26936 20594 26988
rect 20625 26979 20683 26985
rect 20625 26945 20637 26979
rect 20671 26976 20683 26979
rect 21174 26976 21180 26988
rect 20671 26948 21180 26976
rect 20671 26945 20683 26948
rect 20625 26939 20683 26945
rect 21174 26936 21180 26948
rect 21232 26936 21238 26988
rect 22094 26936 22100 26988
rect 22152 26976 22158 26988
rect 25510 26979 25568 26985
rect 25510 26976 25522 26979
rect 22152 26948 22197 26976
rect 23768 26948 25522 26976
rect 22152 26936 22158 26948
rect 19334 26908 19340 26920
rect 19076 26880 19340 26908
rect 17451 26877 17463 26880
rect 17405 26871 17463 26877
rect 19334 26868 19340 26880
rect 19392 26868 19398 26920
rect 21913 26911 21971 26917
rect 21913 26877 21925 26911
rect 21959 26908 21971 26911
rect 22186 26908 22192 26920
rect 21959 26880 22192 26908
rect 21959 26877 21971 26880
rect 21913 26871 21971 26877
rect 22186 26868 22192 26880
rect 22244 26908 22250 26920
rect 22830 26908 22836 26920
rect 22244 26880 22836 26908
rect 22244 26868 22250 26880
rect 22830 26868 22836 26880
rect 22888 26868 22894 26920
rect 10226 26840 10232 26852
rect 10187 26812 10232 26840
rect 10226 26800 10232 26812
rect 10284 26800 10290 26852
rect 11793 26843 11851 26849
rect 11793 26809 11805 26843
rect 11839 26840 11851 26843
rect 23768 26840 23796 26948
rect 25510 26945 25522 26948
rect 25556 26945 25568 26979
rect 25510 26939 25568 26945
rect 27614 26936 27620 26988
rect 27672 26976 27678 26988
rect 28086 26979 28144 26985
rect 28086 26976 28098 26979
rect 27672 26948 28098 26976
rect 27672 26936 27678 26948
rect 28086 26945 28098 26948
rect 28132 26945 28144 26979
rect 28086 26939 28144 26945
rect 28353 26979 28411 26985
rect 28353 26945 28365 26979
rect 28399 26976 28411 26979
rect 29270 26976 29276 26988
rect 28399 26948 29276 26976
rect 28399 26945 28411 26948
rect 28353 26939 28411 26945
rect 29270 26936 29276 26948
rect 29328 26976 29334 26988
rect 29733 26979 29791 26985
rect 29733 26976 29745 26979
rect 29328 26948 29745 26976
rect 29328 26936 29334 26948
rect 29733 26945 29745 26948
rect 29779 26945 29791 26979
rect 33226 26976 33232 26988
rect 33284 26985 33290 26988
rect 33520 26985 33548 27016
rect 33196 26948 33232 26976
rect 29733 26939 29791 26945
rect 33226 26936 33232 26948
rect 33284 26939 33296 26985
rect 33505 26979 33563 26985
rect 33505 26945 33517 26979
rect 33551 26976 33563 26979
rect 33965 26979 34023 26985
rect 33965 26976 33977 26979
rect 33551 26948 33977 26976
rect 33551 26945 33563 26948
rect 33505 26939 33563 26945
rect 33965 26945 33977 26948
rect 34011 26945 34023 26979
rect 33965 26939 34023 26945
rect 33284 26936 33290 26939
rect 34054 26936 34060 26988
rect 34112 26976 34118 26988
rect 34221 26979 34279 26985
rect 34221 26976 34233 26979
rect 34112 26948 34233 26976
rect 34112 26936 34118 26948
rect 34221 26945 34233 26948
rect 34267 26945 34279 26979
rect 34221 26939 34279 26945
rect 25777 26911 25835 26917
rect 25777 26877 25789 26911
rect 25823 26908 25835 26911
rect 26234 26908 26240 26920
rect 25823 26880 26240 26908
rect 25823 26877 25835 26880
rect 25777 26871 25835 26877
rect 26234 26868 26240 26880
rect 26292 26868 26298 26920
rect 26970 26840 26976 26852
rect 11839 26812 23796 26840
rect 26931 26812 26976 26840
rect 11839 26809 11851 26812
rect 11793 26803 11851 26809
rect 26970 26800 26976 26812
rect 27028 26800 27034 26852
rect 8754 26772 8760 26784
rect 8715 26744 8760 26772
rect 8754 26732 8760 26744
rect 8812 26732 8818 26784
rect 14734 26772 14740 26784
rect 14695 26744 14740 26772
rect 14734 26732 14740 26744
rect 14792 26732 14798 26784
rect 15194 26732 15200 26784
rect 15252 26772 15258 26784
rect 15933 26775 15991 26781
rect 15933 26772 15945 26775
rect 15252 26744 15945 26772
rect 15252 26732 15258 26744
rect 15933 26741 15945 26744
rect 15979 26772 15991 26775
rect 16390 26772 16396 26784
rect 15979 26744 16396 26772
rect 15979 26741 15991 26744
rect 15933 26735 15991 26741
rect 16390 26732 16396 26744
rect 16448 26732 16454 26784
rect 16942 26772 16948 26784
rect 16855 26744 16948 26772
rect 16942 26732 16948 26744
rect 17000 26772 17006 26784
rect 17954 26772 17960 26784
rect 17000 26744 17960 26772
rect 17000 26732 17006 26744
rect 17954 26732 17960 26744
rect 18012 26732 18018 26784
rect 18322 26772 18328 26784
rect 18283 26744 18328 26772
rect 18322 26732 18328 26744
rect 18380 26732 18386 26784
rect 19889 26775 19947 26781
rect 19889 26741 19901 26775
rect 19935 26772 19947 26775
rect 22186 26772 22192 26784
rect 19935 26744 22192 26772
rect 19935 26741 19947 26744
rect 19889 26735 19947 26741
rect 22186 26732 22192 26744
rect 22244 26732 22250 26784
rect 22281 26775 22339 26781
rect 22281 26741 22293 26775
rect 22327 26772 22339 26775
rect 22462 26772 22468 26784
rect 22327 26744 22468 26772
rect 22327 26741 22339 26744
rect 22281 26735 22339 26741
rect 22462 26732 22468 26744
rect 22520 26732 22526 26784
rect 22830 26772 22836 26784
rect 22791 26744 22836 26772
rect 22830 26732 22836 26744
rect 22888 26732 22894 26784
rect 23198 26732 23204 26784
rect 23256 26772 23262 26784
rect 24397 26775 24455 26781
rect 24397 26772 24409 26775
rect 23256 26744 24409 26772
rect 23256 26732 23262 26744
rect 24397 26741 24409 26744
rect 24443 26741 24455 26775
rect 24397 26735 24455 26741
rect 30650 26732 30656 26784
rect 30708 26772 30714 26784
rect 31113 26775 31171 26781
rect 31113 26772 31125 26775
rect 30708 26744 31125 26772
rect 30708 26732 30714 26744
rect 31113 26741 31125 26744
rect 31159 26741 31171 26775
rect 31113 26735 31171 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 9122 26568 9128 26580
rect 9083 26540 9128 26568
rect 9122 26528 9128 26540
rect 9180 26528 9186 26580
rect 11238 26568 11244 26580
rect 11199 26540 11244 26568
rect 11238 26528 11244 26540
rect 11296 26528 11302 26580
rect 17126 26568 17132 26580
rect 17087 26540 17132 26568
rect 17126 26528 17132 26540
rect 17184 26528 17190 26580
rect 19058 26528 19064 26580
rect 19116 26568 19122 26580
rect 19116 26540 19564 26568
rect 19116 26528 19122 26540
rect 11882 26500 11888 26512
rect 10336 26472 11100 26500
rect 11843 26472 11888 26500
rect 9582 26392 9588 26444
rect 9640 26432 9646 26444
rect 9677 26435 9735 26441
rect 9677 26432 9689 26435
rect 9640 26404 9689 26432
rect 9640 26392 9646 26404
rect 9677 26401 9689 26404
rect 9723 26401 9735 26435
rect 9677 26395 9735 26401
rect 7374 26324 7380 26376
rect 7432 26364 7438 26376
rect 10336 26373 10364 26472
rect 10873 26435 10931 26441
rect 10873 26401 10885 26435
rect 10919 26432 10931 26435
rect 10962 26432 10968 26444
rect 10919 26404 10968 26432
rect 10919 26401 10931 26404
rect 10873 26395 10931 26401
rect 10962 26392 10968 26404
rect 11020 26392 11026 26444
rect 11072 26432 11100 26472
rect 11882 26460 11888 26472
rect 11940 26460 11946 26512
rect 14921 26503 14979 26509
rect 14921 26469 14933 26503
rect 14967 26500 14979 26503
rect 14967 26472 17908 26500
rect 14967 26469 14979 26472
rect 14921 26463 14979 26469
rect 11072 26404 17816 26432
rect 9493 26367 9551 26373
rect 9493 26364 9505 26367
rect 7432 26336 9505 26364
rect 7432 26324 7438 26336
rect 9493 26333 9505 26336
rect 9539 26364 9551 26367
rect 10321 26367 10379 26373
rect 10321 26364 10333 26367
rect 9539 26336 10333 26364
rect 9539 26333 9551 26336
rect 9493 26327 9551 26333
rect 10321 26333 10333 26336
rect 10367 26333 10379 26367
rect 10321 26327 10379 26333
rect 11057 26367 11115 26373
rect 11057 26333 11069 26367
rect 11103 26364 11115 26367
rect 11514 26364 11520 26376
rect 11103 26336 11520 26364
rect 11103 26333 11115 26336
rect 11057 26327 11115 26333
rect 11514 26324 11520 26336
rect 11572 26324 11578 26376
rect 11698 26364 11704 26376
rect 11659 26336 11704 26364
rect 11698 26324 11704 26336
rect 11756 26324 11762 26376
rect 12250 26324 12256 26376
rect 12308 26364 12314 26376
rect 12894 26364 12900 26376
rect 12308 26336 12900 26364
rect 12308 26324 12314 26336
rect 12894 26324 12900 26336
rect 12952 26324 12958 26376
rect 14734 26364 14740 26376
rect 14695 26336 14740 26364
rect 14734 26324 14740 26336
rect 14792 26324 14798 26376
rect 16482 26324 16488 26376
rect 16540 26364 16546 26376
rect 16761 26367 16819 26373
rect 16761 26364 16773 26367
rect 16540 26336 16773 26364
rect 16540 26324 16546 26336
rect 16761 26333 16773 26336
rect 16807 26333 16819 26367
rect 16942 26364 16948 26376
rect 16903 26336 16948 26364
rect 16761 26327 16819 26333
rect 16942 26324 16948 26336
rect 17000 26324 17006 26376
rect 9585 26299 9643 26305
rect 9585 26265 9597 26299
rect 9631 26296 9643 26299
rect 9858 26296 9864 26308
rect 9631 26268 9864 26296
rect 9631 26265 9643 26268
rect 9585 26259 9643 26265
rect 9858 26256 9864 26268
rect 9916 26256 9922 26308
rect 12912 26228 12940 26324
rect 13170 26296 13176 26308
rect 13131 26268 13176 26296
rect 13170 26256 13176 26268
rect 13228 26256 13234 26308
rect 16301 26299 16359 26305
rect 16301 26265 16313 26299
rect 16347 26296 16359 26299
rect 17126 26296 17132 26308
rect 16347 26268 17132 26296
rect 16347 26265 16359 26268
rect 16301 26259 16359 26265
rect 17126 26256 17132 26268
rect 17184 26256 17190 26308
rect 13814 26228 13820 26240
rect 12912 26200 13820 26228
rect 13814 26188 13820 26200
rect 13872 26188 13878 26240
rect 17788 26228 17816 26404
rect 17880 26296 17908 26472
rect 18506 26460 18512 26512
rect 18564 26500 18570 26512
rect 18601 26503 18659 26509
rect 18601 26500 18613 26503
rect 18564 26472 18613 26500
rect 18564 26460 18570 26472
rect 18601 26469 18613 26472
rect 18647 26469 18659 26503
rect 19536 26500 19564 26540
rect 19610 26528 19616 26580
rect 19668 26568 19674 26580
rect 19978 26568 19984 26580
rect 19668 26540 19984 26568
rect 19668 26528 19674 26540
rect 19978 26528 19984 26540
rect 20036 26568 20042 26580
rect 20438 26568 20444 26580
rect 20036 26540 20444 26568
rect 20036 26528 20042 26540
rect 20438 26528 20444 26540
rect 20496 26528 20502 26580
rect 21174 26568 21180 26580
rect 21135 26540 21180 26568
rect 21174 26528 21180 26540
rect 21232 26528 21238 26580
rect 22186 26528 22192 26580
rect 22244 26568 22250 26580
rect 28994 26568 29000 26580
rect 22244 26540 29000 26568
rect 22244 26528 22250 26540
rect 28994 26528 29000 26540
rect 29052 26528 29058 26580
rect 36630 26528 36636 26580
rect 36688 26568 36694 26580
rect 36998 26568 37004 26580
rect 36688 26540 37004 26568
rect 36688 26528 36694 26540
rect 36998 26528 37004 26540
rect 37056 26568 37062 26580
rect 37645 26571 37703 26577
rect 37645 26568 37657 26571
rect 37056 26540 37657 26568
rect 37056 26528 37062 26540
rect 37645 26537 37657 26540
rect 37691 26537 37703 26571
rect 37645 26531 37703 26537
rect 23750 26500 23756 26512
rect 19536 26472 23756 26500
rect 18601 26463 18659 26469
rect 23750 26460 23756 26472
rect 23808 26460 23814 26512
rect 33226 26460 33232 26512
rect 33284 26500 33290 26512
rect 33410 26500 33416 26512
rect 33284 26472 33416 26500
rect 33284 26460 33290 26472
rect 33410 26460 33416 26472
rect 33468 26460 33474 26512
rect 17954 26392 17960 26444
rect 18012 26432 18018 26444
rect 19429 26435 19487 26441
rect 19429 26432 19441 26435
rect 18012 26404 19441 26432
rect 18012 26392 18018 26404
rect 19429 26401 19441 26404
rect 19475 26432 19487 26435
rect 19518 26432 19524 26444
rect 19475 26404 19524 26432
rect 19475 26401 19487 26404
rect 19429 26395 19487 26401
rect 19518 26392 19524 26404
rect 19576 26392 19582 26444
rect 20162 26392 20168 26444
rect 20220 26432 20226 26444
rect 21729 26435 21787 26441
rect 21729 26432 21741 26435
rect 20220 26404 21741 26432
rect 20220 26392 20226 26404
rect 21729 26401 21741 26404
rect 21775 26401 21787 26435
rect 21729 26395 21787 26401
rect 24302 26392 24308 26444
rect 24360 26432 24366 26444
rect 31938 26432 31944 26444
rect 24360 26404 31944 26432
rect 24360 26392 24366 26404
rect 31938 26392 31944 26404
rect 31996 26392 32002 26444
rect 32306 26392 32312 26444
rect 32364 26432 32370 26444
rect 32953 26435 33011 26441
rect 32953 26432 32965 26435
rect 32364 26404 32965 26432
rect 32364 26392 32370 26404
rect 32953 26401 32965 26404
rect 32999 26432 33011 26435
rect 33042 26432 33048 26444
rect 32999 26404 33048 26432
rect 32999 26401 33011 26404
rect 32953 26395 33011 26401
rect 33042 26392 33048 26404
rect 33100 26392 33106 26444
rect 18233 26367 18291 26373
rect 18233 26333 18245 26367
rect 18279 26364 18291 26367
rect 19242 26364 19248 26376
rect 18279 26336 19248 26364
rect 18279 26333 18291 26336
rect 18233 26327 18291 26333
rect 19242 26324 19248 26336
rect 19300 26364 19306 26376
rect 20346 26364 20352 26376
rect 19300 26336 20352 26364
rect 19300 26324 19306 26336
rect 20346 26324 20352 26336
rect 20404 26324 20410 26376
rect 21450 26324 21456 26376
rect 21508 26364 21514 26376
rect 21545 26367 21603 26373
rect 21545 26364 21557 26367
rect 21508 26336 21557 26364
rect 21508 26324 21514 26336
rect 21545 26333 21557 26336
rect 21591 26364 21603 26367
rect 27798 26364 27804 26376
rect 21591 26336 23060 26364
rect 27759 26336 27804 26364
rect 21591 26333 21603 26336
rect 21545 26327 21603 26333
rect 23032 26308 23060 26336
rect 27798 26324 27804 26336
rect 27856 26364 27862 26376
rect 30374 26364 30380 26376
rect 27856 26336 30380 26364
rect 27856 26324 27862 26336
rect 30374 26324 30380 26336
rect 30432 26364 30438 26376
rect 31205 26367 31263 26373
rect 31205 26364 31217 26367
rect 30432 26336 31217 26364
rect 30432 26324 30438 26336
rect 31205 26333 31217 26336
rect 31251 26333 31263 26367
rect 31205 26327 31263 26333
rect 18141 26299 18199 26305
rect 17880 26268 18092 26296
rect 17954 26228 17960 26240
rect 17788 26200 17960 26228
rect 17954 26188 17960 26200
rect 18012 26188 18018 26240
rect 18064 26228 18092 26268
rect 18141 26265 18153 26299
rect 18187 26296 18199 26299
rect 18322 26296 18328 26308
rect 18187 26268 18328 26296
rect 18187 26265 18199 26268
rect 18141 26259 18199 26265
rect 18322 26256 18328 26268
rect 18380 26256 18386 26308
rect 19058 26296 19064 26308
rect 18432 26268 19064 26296
rect 18432 26228 18460 26268
rect 19058 26256 19064 26268
rect 19116 26256 19122 26308
rect 19521 26299 19579 26305
rect 19521 26265 19533 26299
rect 19567 26296 19579 26299
rect 20070 26296 20076 26308
rect 19567 26268 20076 26296
rect 19567 26265 19579 26268
rect 19521 26259 19579 26265
rect 20070 26256 20076 26268
rect 20128 26256 20134 26308
rect 21637 26299 21695 26305
rect 21637 26265 21649 26299
rect 21683 26296 21695 26299
rect 22370 26296 22376 26308
rect 21683 26268 22376 26296
rect 21683 26265 21695 26268
rect 21637 26259 21695 26265
rect 22370 26256 22376 26268
rect 22428 26256 22434 26308
rect 23014 26296 23020 26308
rect 22975 26268 23020 26296
rect 23014 26256 23020 26268
rect 23072 26256 23078 26308
rect 26234 26296 26240 26308
rect 26195 26268 26240 26296
rect 26234 26256 26240 26268
rect 26292 26256 26298 26308
rect 31220 26296 31248 26327
rect 31478 26324 31484 26376
rect 31536 26364 31542 26376
rect 33410 26364 33416 26376
rect 31536 26336 33416 26364
rect 31536 26324 31542 26336
rect 33410 26324 33416 26336
rect 33468 26324 33474 26376
rect 35342 26364 35348 26376
rect 35303 26336 35348 26364
rect 35342 26324 35348 26336
rect 35400 26324 35406 26376
rect 33134 26296 33140 26308
rect 31220 26268 33140 26296
rect 33134 26256 33140 26268
rect 33192 26296 33198 26308
rect 36357 26299 36415 26305
rect 36357 26296 36369 26299
rect 33192 26268 36369 26296
rect 33192 26256 33198 26268
rect 36357 26265 36369 26268
rect 36403 26265 36415 26299
rect 36357 26259 36415 26265
rect 19610 26228 19616 26240
rect 18064 26200 18460 26228
rect 19571 26200 19616 26228
rect 19610 26188 19616 26200
rect 19668 26188 19674 26240
rect 19978 26228 19984 26240
rect 19939 26200 19984 26228
rect 19978 26188 19984 26200
rect 20036 26188 20042 26240
rect 35526 26228 35532 26240
rect 35487 26200 35532 26228
rect 35526 26188 35532 26200
rect 35584 26188 35590 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 9309 26027 9367 26033
rect 9309 25993 9321 26027
rect 9355 26024 9367 26027
rect 9490 26024 9496 26036
rect 9355 25996 9496 26024
rect 9355 25993 9367 25996
rect 9309 25987 9367 25993
rect 9490 25984 9496 25996
rect 9548 25984 9554 26036
rect 15838 25984 15844 26036
rect 15896 26024 15902 26036
rect 16025 26027 16083 26033
rect 16025 26024 16037 26027
rect 15896 25996 16037 26024
rect 15896 25984 15902 25996
rect 16025 25993 16037 25996
rect 16071 25993 16083 26027
rect 16025 25987 16083 25993
rect 16669 26027 16727 26033
rect 16669 25993 16681 26027
rect 16715 26024 16727 26027
rect 16942 26024 16948 26036
rect 16715 25996 16948 26024
rect 16715 25993 16727 25996
rect 16669 25987 16727 25993
rect 16040 25956 16068 25987
rect 16942 25984 16948 25996
rect 17000 25984 17006 26036
rect 18325 26027 18383 26033
rect 18325 25993 18337 26027
rect 18371 26024 18383 26027
rect 18414 26024 18420 26036
rect 18371 25996 18420 26024
rect 18371 25993 18383 25996
rect 18325 25987 18383 25993
rect 18414 25984 18420 25996
rect 18472 25984 18478 26036
rect 19058 25984 19064 26036
rect 19116 26024 19122 26036
rect 20530 26024 20536 26036
rect 19116 25996 20536 26024
rect 19116 25984 19122 25996
rect 20530 25984 20536 25996
rect 20588 25984 20594 26036
rect 29089 26027 29147 26033
rect 29089 25993 29101 26027
rect 29135 26024 29147 26027
rect 29270 26024 29276 26036
rect 29135 25996 29276 26024
rect 29135 25993 29147 25996
rect 29089 25987 29147 25993
rect 29270 25984 29276 25996
rect 29328 25984 29334 26036
rect 32125 26027 32183 26033
rect 32125 26024 32137 26027
rect 29380 25996 32137 26024
rect 17034 25956 17040 25968
rect 16040 25928 17040 25956
rect 17034 25916 17040 25928
rect 17092 25916 17098 25968
rect 23014 25916 23020 25968
rect 23072 25956 23078 25968
rect 29380 25956 29408 25996
rect 32125 25993 32137 25996
rect 32171 25993 32183 26027
rect 32125 25987 32183 25993
rect 35526 25984 35532 26036
rect 35584 26024 35590 26036
rect 36722 26024 36728 26036
rect 35584 25996 35664 26024
rect 36683 25996 36728 26024
rect 35584 25984 35590 25996
rect 30374 25956 30380 25968
rect 23072 25928 29408 25956
rect 30335 25928 30380 25956
rect 23072 25916 23078 25928
rect 30374 25916 30380 25928
rect 30432 25916 30438 25968
rect 32306 25916 32312 25968
rect 32364 25956 32370 25968
rect 35636 25965 35664 25996
rect 36722 25984 36728 25996
rect 36780 25984 36786 26036
rect 37826 26024 37832 26036
rect 37787 25996 37832 26024
rect 37826 25984 37832 25996
rect 37884 25984 37890 26036
rect 35612 25959 35670 25965
rect 32364 25928 33548 25956
rect 32364 25916 32370 25928
rect 8754 25848 8760 25900
rect 8812 25888 8818 25900
rect 9125 25891 9183 25897
rect 9125 25888 9137 25891
rect 8812 25860 9137 25888
rect 8812 25848 8818 25860
rect 9125 25857 9137 25860
rect 9171 25857 9183 25891
rect 9125 25851 9183 25857
rect 17402 25848 17408 25900
rect 17460 25888 17466 25900
rect 20717 25891 20775 25897
rect 20717 25888 20729 25891
rect 17460 25860 20729 25888
rect 17460 25848 17466 25860
rect 20717 25857 20729 25860
rect 20763 25888 20775 25891
rect 22189 25891 22247 25897
rect 20763 25860 21864 25888
rect 20763 25857 20775 25860
rect 20717 25851 20775 25857
rect 17126 25820 17132 25832
rect 17087 25792 17132 25820
rect 17126 25780 17132 25792
rect 17184 25780 17190 25832
rect 17221 25823 17279 25829
rect 17221 25789 17233 25823
rect 17267 25789 17279 25823
rect 17221 25783 17279 25789
rect 16482 25712 16488 25764
rect 16540 25752 16546 25764
rect 17236 25752 17264 25783
rect 17954 25780 17960 25832
rect 18012 25820 18018 25832
rect 21836 25829 21864 25860
rect 22189 25857 22201 25891
rect 22235 25888 22247 25891
rect 24946 25888 24952 25900
rect 22235 25860 24952 25888
rect 22235 25857 22247 25860
rect 22189 25851 22247 25857
rect 24946 25848 24952 25860
rect 25004 25848 25010 25900
rect 25222 25848 25228 25900
rect 25280 25897 25286 25900
rect 25280 25888 25292 25897
rect 33249 25891 33307 25897
rect 25280 25860 25325 25888
rect 25280 25851 25292 25860
rect 33249 25857 33261 25891
rect 33295 25888 33307 25891
rect 33410 25888 33416 25900
rect 33295 25860 33416 25888
rect 33295 25857 33307 25860
rect 33249 25851 33307 25857
rect 25280 25848 25286 25851
rect 33410 25848 33416 25860
rect 33468 25848 33474 25900
rect 33520 25897 33548 25928
rect 35612 25925 35624 25959
rect 35658 25925 35670 25959
rect 35612 25919 35670 25925
rect 33505 25891 33563 25897
rect 33505 25857 33517 25891
rect 33551 25857 33563 25891
rect 38010 25888 38016 25900
rect 37971 25860 38016 25888
rect 33505 25851 33563 25857
rect 38010 25848 38016 25860
rect 38068 25848 38074 25900
rect 21821 25823 21879 25829
rect 18012 25792 20668 25820
rect 18012 25780 18018 25792
rect 16540 25724 17264 25752
rect 19889 25755 19947 25761
rect 16540 25712 16546 25724
rect 19889 25721 19901 25755
rect 19935 25752 19947 25755
rect 20070 25752 20076 25764
rect 19935 25724 20076 25752
rect 19935 25721 19947 25724
rect 19889 25715 19947 25721
rect 20070 25712 20076 25724
rect 20128 25752 20134 25764
rect 20530 25752 20536 25764
rect 20128 25724 20536 25752
rect 20128 25712 20134 25724
rect 20530 25712 20536 25724
rect 20588 25712 20594 25764
rect 20640 25752 20668 25792
rect 21821 25789 21833 25823
rect 21867 25789 21879 25823
rect 21821 25783 21879 25789
rect 22281 25823 22339 25829
rect 22281 25789 22293 25823
rect 22327 25820 22339 25823
rect 22554 25820 22560 25832
rect 22327 25792 22560 25820
rect 22327 25789 22339 25792
rect 22281 25783 22339 25789
rect 22554 25780 22560 25792
rect 22612 25780 22618 25832
rect 25501 25823 25559 25829
rect 25501 25789 25513 25823
rect 25547 25820 25559 25823
rect 26234 25820 26240 25832
rect 25547 25792 26240 25820
rect 25547 25789 25559 25792
rect 25501 25783 25559 25789
rect 26234 25780 26240 25792
rect 26292 25780 26298 25832
rect 35345 25823 35403 25829
rect 35345 25789 35357 25823
rect 35391 25789 35403 25823
rect 35345 25783 35403 25789
rect 24121 25755 24179 25761
rect 24121 25752 24133 25755
rect 20640 25724 24133 25752
rect 24121 25721 24133 25724
rect 24167 25721 24179 25755
rect 24121 25715 24179 25721
rect 9858 25644 9864 25696
rect 9916 25684 9922 25696
rect 10137 25687 10195 25693
rect 10137 25684 10149 25687
rect 9916 25656 10149 25684
rect 9916 25644 9922 25656
rect 10137 25653 10149 25656
rect 10183 25653 10195 25687
rect 10778 25684 10784 25696
rect 10691 25656 10784 25684
rect 10137 25647 10195 25653
rect 10778 25644 10784 25656
rect 10836 25684 10842 25696
rect 12158 25684 12164 25696
rect 10836 25656 12164 25684
rect 10836 25644 10842 25656
rect 12158 25644 12164 25656
rect 12216 25644 12222 25696
rect 12342 25644 12348 25696
rect 12400 25684 12406 25696
rect 12437 25687 12495 25693
rect 12437 25684 12449 25687
rect 12400 25656 12449 25684
rect 12400 25644 12406 25656
rect 12437 25653 12449 25656
rect 12483 25653 12495 25687
rect 15562 25684 15568 25696
rect 15523 25656 15568 25684
rect 12437 25647 12495 25653
rect 15562 25644 15568 25656
rect 15620 25644 15626 25696
rect 18877 25687 18935 25693
rect 18877 25653 18889 25687
rect 18923 25684 18935 25687
rect 19058 25684 19064 25696
rect 18923 25656 19064 25684
rect 18923 25653 18935 25656
rect 18877 25647 18935 25653
rect 19058 25644 19064 25656
rect 19116 25644 19122 25696
rect 20162 25644 20168 25696
rect 20220 25684 20226 25696
rect 20441 25687 20499 25693
rect 20441 25684 20453 25687
rect 20220 25656 20453 25684
rect 20220 25644 20226 25656
rect 20441 25653 20453 25656
rect 20487 25653 20499 25687
rect 20441 25647 20499 25653
rect 34606 25644 34612 25696
rect 34664 25684 34670 25696
rect 34790 25684 34796 25696
rect 34664 25656 34796 25684
rect 34664 25644 34670 25656
rect 34790 25644 34796 25656
rect 34848 25644 34854 25696
rect 35360 25684 35388 25783
rect 36354 25684 36360 25696
rect 35360 25656 36360 25684
rect 36354 25644 36360 25656
rect 36412 25684 36418 25696
rect 36630 25684 36636 25696
rect 36412 25656 36636 25684
rect 36412 25644 36418 25656
rect 36630 25644 36636 25656
rect 36688 25644 36694 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 8570 25440 8576 25492
rect 8628 25480 8634 25492
rect 8941 25483 8999 25489
rect 8941 25480 8953 25483
rect 8628 25452 8953 25480
rect 8628 25440 8634 25452
rect 8941 25449 8953 25452
rect 8987 25449 8999 25483
rect 8941 25443 8999 25449
rect 11054 25440 11060 25492
rect 11112 25480 11118 25492
rect 11609 25483 11667 25489
rect 11609 25480 11621 25483
rect 11112 25452 11621 25480
rect 11112 25440 11118 25452
rect 11609 25449 11621 25452
rect 11655 25449 11667 25483
rect 12897 25483 12955 25489
rect 12897 25480 12909 25483
rect 11609 25443 11667 25449
rect 12406 25452 12909 25480
rect 10226 25412 10232 25424
rect 9324 25384 10232 25412
rect 8938 25304 8944 25356
rect 8996 25344 9002 25356
rect 9324 25344 9352 25384
rect 10226 25372 10232 25384
rect 10284 25372 10290 25424
rect 12158 25372 12164 25424
rect 12216 25412 12222 25424
rect 12406 25412 12434 25452
rect 12897 25449 12909 25452
rect 12943 25480 12955 25483
rect 13722 25480 13728 25492
rect 12943 25452 13728 25480
rect 12943 25449 12955 25452
rect 12897 25443 12955 25449
rect 13722 25440 13728 25452
rect 13780 25440 13786 25492
rect 15470 25440 15476 25492
rect 15528 25480 15534 25492
rect 15841 25483 15899 25489
rect 15841 25480 15853 25483
rect 15528 25452 15853 25480
rect 15528 25440 15534 25452
rect 15841 25449 15853 25452
rect 15887 25449 15899 25483
rect 15841 25443 15899 25449
rect 18693 25483 18751 25489
rect 18693 25449 18705 25483
rect 18739 25480 18751 25483
rect 18966 25480 18972 25492
rect 18739 25452 18972 25480
rect 18739 25449 18751 25452
rect 18693 25443 18751 25449
rect 18966 25440 18972 25452
rect 19024 25440 19030 25492
rect 26237 25483 26295 25489
rect 26237 25480 26249 25483
rect 22066 25452 26249 25480
rect 13446 25412 13452 25424
rect 12216 25384 12434 25412
rect 13407 25384 13452 25412
rect 12216 25372 12222 25384
rect 13446 25372 13452 25384
rect 13504 25372 13510 25424
rect 20162 25412 20168 25424
rect 18064 25384 20168 25412
rect 9582 25344 9588 25356
rect 8996 25316 9352 25344
rect 9543 25316 9588 25344
rect 8996 25304 9002 25316
rect 9324 25285 9352 25316
rect 9582 25304 9588 25316
rect 9640 25304 9646 25356
rect 12250 25344 12256 25356
rect 12211 25316 12256 25344
rect 12250 25304 12256 25316
rect 12308 25304 12314 25356
rect 12434 25304 12440 25356
rect 12492 25344 12498 25356
rect 12492 25316 14964 25344
rect 12492 25304 12498 25316
rect 9309 25279 9367 25285
rect 9309 25245 9321 25279
rect 9355 25245 9367 25279
rect 9309 25239 9367 25245
rect 11977 25279 12035 25285
rect 11977 25245 11989 25279
rect 12023 25276 12035 25279
rect 13446 25276 13452 25288
rect 12023 25248 13452 25276
rect 12023 25245 12035 25248
rect 11977 25239 12035 25245
rect 13446 25236 13452 25248
rect 13504 25236 13510 25288
rect 14936 25276 14964 25316
rect 15010 25304 15016 25356
rect 15068 25344 15074 25356
rect 15197 25347 15255 25353
rect 15197 25344 15209 25347
rect 15068 25316 15209 25344
rect 15068 25304 15074 25316
rect 15197 25313 15209 25316
rect 15243 25344 15255 25347
rect 16482 25344 16488 25356
rect 15243 25316 16488 25344
rect 15243 25313 15255 25316
rect 15197 25307 15255 25313
rect 16482 25304 16488 25316
rect 16540 25344 16546 25356
rect 17129 25347 17187 25353
rect 17129 25344 17141 25347
rect 16540 25316 17141 25344
rect 16540 25304 16546 25316
rect 17129 25313 17141 25316
rect 17175 25313 17187 25347
rect 17129 25307 17187 25313
rect 17954 25304 17960 25356
rect 18012 25344 18018 25356
rect 18064 25353 18092 25384
rect 20162 25372 20168 25384
rect 20220 25372 20226 25424
rect 20346 25372 20352 25424
rect 20404 25412 20410 25424
rect 22066 25412 22094 25452
rect 26237 25449 26249 25452
rect 26283 25449 26295 25483
rect 26237 25443 26295 25449
rect 33873 25483 33931 25489
rect 33873 25449 33885 25483
rect 33919 25480 33931 25483
rect 34054 25480 34060 25492
rect 33919 25452 34060 25480
rect 33919 25449 33931 25452
rect 33873 25443 33931 25449
rect 34054 25440 34060 25452
rect 34112 25440 34118 25492
rect 35342 25480 35348 25492
rect 35303 25452 35348 25480
rect 35342 25440 35348 25452
rect 35400 25440 35406 25492
rect 22646 25412 22652 25424
rect 20404 25384 22094 25412
rect 22607 25384 22652 25412
rect 20404 25372 20410 25384
rect 22646 25372 22652 25384
rect 22704 25372 22710 25424
rect 24397 25415 24455 25421
rect 24397 25381 24409 25415
rect 24443 25381 24455 25415
rect 24397 25375 24455 25381
rect 34885 25415 34943 25421
rect 34885 25381 34897 25415
rect 34931 25412 34943 25415
rect 35710 25412 35716 25424
rect 34931 25384 35716 25412
rect 34931 25381 34943 25384
rect 34885 25375 34943 25381
rect 18049 25347 18107 25353
rect 18049 25344 18061 25347
rect 18012 25316 18061 25344
rect 18012 25304 18018 25316
rect 18049 25313 18061 25316
rect 18095 25313 18107 25347
rect 18049 25307 18107 25313
rect 18138 25304 18144 25356
rect 18196 25344 18202 25356
rect 24412 25344 24440 25375
rect 35710 25372 35716 25384
rect 35768 25372 35774 25424
rect 18196 25316 24440 25344
rect 18196 25304 18202 25316
rect 29270 25304 29276 25356
rect 29328 25344 29334 25356
rect 29549 25347 29607 25353
rect 29549 25344 29561 25347
rect 29328 25316 29561 25344
rect 29328 25304 29334 25316
rect 29549 25313 29561 25316
rect 29595 25313 29607 25347
rect 29549 25307 29607 25313
rect 36354 25304 36360 25356
rect 36412 25344 36418 25356
rect 36725 25347 36783 25353
rect 36725 25344 36737 25347
rect 36412 25316 36737 25344
rect 36412 25304 36418 25316
rect 36725 25313 36737 25316
rect 36771 25313 36783 25347
rect 36725 25307 36783 25313
rect 15473 25279 15531 25285
rect 15473 25276 15485 25279
rect 14936 25248 15485 25276
rect 15473 25245 15485 25248
rect 15519 25276 15531 25279
rect 16666 25276 16672 25288
rect 15519 25248 16672 25276
rect 15519 25245 15531 25248
rect 15473 25239 15531 25245
rect 16666 25236 16672 25248
rect 16724 25236 16730 25288
rect 17402 25276 17408 25288
rect 17363 25248 17408 25276
rect 17402 25236 17408 25248
rect 17460 25236 17466 25288
rect 18325 25279 18383 25285
rect 18325 25245 18337 25279
rect 18371 25276 18383 25279
rect 18414 25276 18420 25288
rect 18371 25248 18420 25276
rect 18371 25245 18383 25248
rect 18325 25239 18383 25245
rect 18414 25236 18420 25248
rect 18472 25236 18478 25288
rect 20622 25276 20628 25288
rect 20364 25248 20628 25276
rect 9401 25211 9459 25217
rect 9401 25177 9413 25211
rect 9447 25208 9459 25211
rect 15381 25211 15439 25217
rect 9447 25180 10456 25208
rect 9447 25177 9459 25180
rect 9401 25171 9459 25177
rect 10428 25152 10456 25180
rect 15381 25177 15393 25211
rect 15427 25208 15439 25211
rect 15562 25208 15568 25220
rect 15427 25180 15568 25208
rect 15427 25177 15439 25180
rect 15381 25171 15439 25177
rect 15562 25168 15568 25180
rect 15620 25208 15626 25220
rect 16298 25208 16304 25220
rect 15620 25180 16304 25208
rect 15620 25168 15626 25180
rect 16298 25168 16304 25180
rect 16356 25168 16362 25220
rect 16577 25211 16635 25217
rect 16577 25177 16589 25211
rect 16623 25208 16635 25211
rect 19521 25211 19579 25217
rect 16623 25180 18092 25208
rect 16623 25177 16635 25180
rect 16577 25171 16635 25177
rect 18064 25152 18092 25180
rect 19521 25177 19533 25211
rect 19567 25208 19579 25211
rect 20070 25208 20076 25220
rect 19567 25180 20076 25208
rect 19567 25177 19579 25180
rect 19521 25171 19579 25177
rect 20070 25168 20076 25180
rect 20128 25168 20134 25220
rect 20364 25152 20392 25248
rect 20622 25236 20628 25248
rect 20680 25236 20686 25288
rect 22462 25276 22468 25288
rect 22423 25248 22468 25276
rect 22462 25236 22468 25248
rect 22520 25236 22526 25288
rect 23750 25236 23756 25288
rect 23808 25276 23814 25288
rect 25510 25279 25568 25285
rect 25510 25276 25522 25279
rect 23808 25248 25522 25276
rect 23808 25236 23814 25248
rect 25510 25245 25522 25248
rect 25556 25245 25568 25279
rect 25510 25239 25568 25245
rect 25777 25279 25835 25285
rect 25777 25245 25789 25279
rect 25823 25276 25835 25279
rect 26234 25276 26240 25288
rect 25823 25248 26240 25276
rect 25823 25245 25835 25248
rect 25777 25239 25835 25245
rect 26234 25236 26240 25248
rect 26292 25276 26298 25288
rect 27617 25279 27675 25285
rect 27617 25276 27629 25279
rect 26292 25248 27629 25276
rect 26292 25236 26298 25248
rect 27617 25245 27629 25248
rect 27663 25245 27675 25279
rect 27617 25239 27675 25245
rect 28994 25236 29000 25288
rect 29052 25276 29058 25288
rect 29805 25279 29863 25285
rect 29805 25276 29817 25279
rect 29052 25248 29817 25276
rect 29052 25236 29058 25248
rect 29805 25245 29817 25248
rect 29851 25245 29863 25279
rect 32769 25279 32827 25285
rect 32769 25276 32781 25279
rect 29805 25239 29863 25245
rect 32324 25248 32781 25276
rect 32324 25220 32352 25248
rect 32769 25245 32781 25248
rect 32815 25245 32827 25279
rect 33686 25276 33692 25288
rect 33647 25248 33692 25276
rect 32769 25239 32827 25245
rect 33686 25236 33692 25248
rect 33744 25236 33750 25288
rect 34698 25276 34704 25288
rect 34659 25248 34704 25276
rect 34698 25236 34704 25248
rect 34756 25236 34762 25288
rect 35526 25276 35532 25288
rect 35487 25248 35532 25276
rect 35526 25236 35532 25248
rect 35584 25236 35590 25288
rect 35710 25276 35716 25288
rect 35671 25248 35716 25276
rect 35710 25236 35716 25248
rect 35768 25276 35774 25288
rect 36173 25279 36231 25285
rect 36173 25276 36185 25279
rect 35768 25248 36185 25276
rect 35768 25236 35774 25248
rect 36173 25245 36185 25248
rect 36219 25245 36231 25279
rect 36173 25239 36231 25245
rect 22186 25168 22192 25220
rect 22244 25208 22250 25220
rect 22830 25208 22836 25220
rect 22244 25180 22836 25208
rect 22244 25168 22250 25180
rect 22830 25168 22836 25180
rect 22888 25208 22894 25220
rect 23201 25211 23259 25217
rect 23201 25208 23213 25211
rect 22888 25180 23213 25208
rect 22888 25168 22894 25180
rect 23201 25177 23213 25180
rect 23247 25208 23259 25211
rect 24394 25208 24400 25220
rect 23247 25180 24400 25208
rect 23247 25177 23259 25180
rect 23201 25171 23259 25177
rect 24394 25168 24400 25180
rect 24452 25168 24458 25220
rect 26326 25168 26332 25220
rect 26384 25208 26390 25220
rect 27350 25211 27408 25217
rect 27350 25208 27362 25211
rect 26384 25180 27362 25208
rect 26384 25168 26390 25180
rect 27350 25177 27362 25180
rect 27396 25177 27408 25211
rect 27350 25171 27408 25177
rect 32306 25168 32312 25220
rect 32364 25168 32370 25220
rect 32502 25211 32560 25217
rect 32502 25208 32514 25211
rect 32416 25180 32514 25208
rect 10410 25100 10416 25152
rect 10468 25140 10474 25152
rect 10689 25143 10747 25149
rect 10689 25140 10701 25143
rect 10468 25112 10701 25140
rect 10468 25100 10474 25112
rect 10689 25109 10701 25112
rect 10735 25109 10747 25143
rect 10689 25103 10747 25109
rect 12069 25143 12127 25149
rect 12069 25109 12081 25143
rect 12115 25140 12127 25143
rect 12342 25140 12348 25152
rect 12115 25112 12348 25140
rect 12115 25109 12127 25112
rect 12069 25103 12127 25109
rect 12342 25100 12348 25112
rect 12400 25100 12406 25152
rect 14090 25140 14096 25152
rect 14051 25112 14096 25140
rect 14090 25100 14096 25112
rect 14148 25100 14154 25152
rect 18046 25100 18052 25152
rect 18104 25140 18110 25152
rect 18233 25143 18291 25149
rect 18233 25140 18245 25143
rect 18104 25112 18245 25140
rect 18104 25100 18110 25112
rect 18233 25109 18245 25112
rect 18279 25109 18291 25143
rect 18233 25103 18291 25109
rect 19981 25143 20039 25149
rect 19981 25109 19993 25143
rect 20027 25140 20039 25143
rect 20346 25140 20352 25152
rect 20027 25112 20352 25140
rect 20027 25109 20039 25112
rect 19981 25103 20039 25109
rect 20346 25100 20352 25112
rect 20404 25100 20410 25152
rect 20622 25140 20628 25152
rect 20583 25112 20628 25140
rect 20622 25100 20628 25112
rect 20680 25100 20686 25152
rect 20990 25100 20996 25152
rect 21048 25140 21054 25152
rect 21085 25143 21143 25149
rect 21085 25140 21097 25143
rect 21048 25112 21097 25140
rect 21048 25100 21054 25112
rect 21085 25109 21097 25112
rect 21131 25109 21143 25143
rect 21818 25140 21824 25152
rect 21779 25112 21824 25140
rect 21085 25103 21143 25109
rect 21818 25100 21824 25112
rect 21876 25100 21882 25152
rect 23658 25100 23664 25152
rect 23716 25140 23722 25152
rect 23753 25143 23811 25149
rect 23753 25140 23765 25143
rect 23716 25112 23765 25140
rect 23716 25100 23722 25112
rect 23753 25109 23765 25112
rect 23799 25140 23811 25143
rect 30650 25140 30656 25152
rect 23799 25112 30656 25140
rect 23799 25109 23811 25112
rect 23753 25103 23811 25109
rect 30650 25100 30656 25112
rect 30708 25100 30714 25152
rect 30926 25140 30932 25152
rect 30887 25112 30932 25140
rect 30926 25100 30932 25112
rect 30984 25100 30990 25152
rect 31018 25100 31024 25152
rect 31076 25140 31082 25152
rect 31389 25143 31447 25149
rect 31389 25140 31401 25143
rect 31076 25112 31401 25140
rect 31076 25100 31082 25112
rect 31389 25109 31401 25112
rect 31435 25109 31447 25143
rect 31389 25103 31447 25109
rect 31938 25100 31944 25152
rect 31996 25140 32002 25152
rect 32416 25140 32444 25180
rect 32502 25177 32514 25180
rect 32548 25177 32560 25211
rect 32502 25171 32560 25177
rect 35986 25168 35992 25220
rect 36044 25208 36050 25220
rect 36970 25211 37028 25217
rect 36970 25208 36982 25211
rect 36044 25180 36982 25208
rect 36044 25168 36050 25180
rect 36970 25177 36982 25180
rect 37016 25177 37028 25211
rect 36970 25171 37028 25177
rect 31996 25112 32444 25140
rect 31996 25100 32002 25112
rect 37826 25100 37832 25152
rect 37884 25140 37890 25152
rect 38105 25143 38163 25149
rect 38105 25140 38117 25143
rect 37884 25112 38117 25140
rect 37884 25100 37890 25112
rect 38105 25109 38117 25112
rect 38151 25140 38163 25143
rect 38194 25140 38200 25152
rect 38151 25112 38200 25140
rect 38151 25109 38163 25112
rect 38105 25103 38163 25109
rect 38194 25100 38200 25112
rect 38252 25100 38258 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 9582 24896 9588 24948
rect 9640 24936 9646 24948
rect 9861 24939 9919 24945
rect 9861 24936 9873 24939
rect 9640 24908 9873 24936
rect 9640 24896 9646 24908
rect 9861 24905 9873 24908
rect 9907 24936 9919 24939
rect 10778 24936 10784 24948
rect 9907 24908 10784 24936
rect 9907 24905 9919 24908
rect 9861 24899 9919 24905
rect 10778 24896 10784 24908
rect 10836 24896 10842 24948
rect 13630 24936 13636 24948
rect 13591 24908 13636 24936
rect 13630 24896 13636 24908
rect 13688 24896 13694 24948
rect 14826 24936 14832 24948
rect 14787 24908 14832 24936
rect 14826 24896 14832 24908
rect 14884 24936 14890 24948
rect 15657 24939 15715 24945
rect 15657 24936 15669 24939
rect 14884 24908 15669 24936
rect 14884 24896 14890 24908
rect 15657 24905 15669 24908
rect 15703 24905 15715 24939
rect 15657 24899 15715 24905
rect 17494 24896 17500 24948
rect 17552 24936 17558 24948
rect 20441 24939 20499 24945
rect 20441 24936 20453 24939
rect 17552 24908 20453 24936
rect 17552 24896 17558 24908
rect 20441 24905 20453 24908
rect 20487 24936 20499 24939
rect 20990 24936 20996 24948
rect 20487 24908 20996 24936
rect 20487 24905 20499 24908
rect 20441 24899 20499 24905
rect 20990 24896 20996 24908
rect 21048 24936 21054 24948
rect 31018 24936 31024 24948
rect 21048 24908 31024 24936
rect 21048 24896 21054 24908
rect 31018 24896 31024 24908
rect 31076 24896 31082 24948
rect 37642 24896 37648 24948
rect 37700 24936 37706 24948
rect 37737 24939 37795 24945
rect 37737 24936 37749 24939
rect 37700 24908 37749 24936
rect 37700 24896 37706 24908
rect 37737 24905 37749 24908
rect 37783 24905 37795 24939
rect 37737 24899 37795 24905
rect 11422 24828 11428 24880
rect 11480 24868 11486 24880
rect 11885 24871 11943 24877
rect 11885 24868 11897 24871
rect 11480 24840 11897 24868
rect 11480 24828 11486 24840
rect 11885 24837 11897 24840
rect 11931 24837 11943 24871
rect 11885 24831 11943 24837
rect 17589 24871 17647 24877
rect 17589 24837 17601 24871
rect 17635 24868 17647 24871
rect 17678 24868 17684 24880
rect 17635 24840 17684 24868
rect 17635 24837 17647 24840
rect 17589 24831 17647 24837
rect 11900 24800 11928 24831
rect 17678 24828 17684 24840
rect 17736 24828 17742 24880
rect 14090 24800 14096 24812
rect 11900 24772 12848 24800
rect 11974 24732 11980 24744
rect 11935 24704 11980 24732
rect 11974 24692 11980 24704
rect 12032 24692 12038 24744
rect 12158 24732 12164 24744
rect 12119 24704 12164 24732
rect 12158 24692 12164 24704
rect 12216 24692 12222 24744
rect 11514 24664 11520 24676
rect 11475 24636 11520 24664
rect 11514 24624 11520 24636
rect 11572 24624 11578 24676
rect 12820 24605 12848 24772
rect 13740 24772 14096 24800
rect 13446 24692 13452 24744
rect 13504 24732 13510 24744
rect 13740 24741 13768 24772
rect 14090 24760 14096 24772
rect 14148 24760 14154 24812
rect 14921 24803 14979 24809
rect 14921 24769 14933 24803
rect 14967 24800 14979 24803
rect 15286 24800 15292 24812
rect 14967 24772 15292 24800
rect 14967 24769 14979 24772
rect 14921 24763 14979 24769
rect 15286 24760 15292 24772
rect 15344 24760 15350 24812
rect 16666 24800 16672 24812
rect 16627 24772 16672 24800
rect 16666 24760 16672 24772
rect 16724 24760 16730 24812
rect 19058 24800 19064 24812
rect 19019 24772 19064 24800
rect 19058 24760 19064 24772
rect 19116 24760 19122 24812
rect 22186 24800 22192 24812
rect 22147 24772 22192 24800
rect 22186 24760 22192 24772
rect 22244 24760 22250 24812
rect 22370 24800 22376 24812
rect 22331 24772 22376 24800
rect 22370 24760 22376 24772
rect 22428 24760 22434 24812
rect 22557 24803 22615 24809
rect 22557 24769 22569 24803
rect 22603 24800 22615 24803
rect 23109 24803 23167 24809
rect 23109 24800 23121 24803
rect 22603 24772 23121 24800
rect 22603 24769 22615 24772
rect 22557 24763 22615 24769
rect 23109 24769 23121 24772
rect 23155 24769 23167 24803
rect 28822 24803 28880 24809
rect 28822 24800 28834 24803
rect 23109 24763 23167 24769
rect 25424 24772 28834 24800
rect 13725 24735 13783 24741
rect 13725 24732 13737 24735
rect 13504 24704 13737 24732
rect 13504 24692 13510 24704
rect 13725 24701 13737 24704
rect 13771 24701 13783 24735
rect 13725 24695 13783 24701
rect 13814 24692 13820 24744
rect 13872 24732 13878 24744
rect 15010 24732 15016 24744
rect 13872 24704 15016 24732
rect 13872 24692 13878 24704
rect 15010 24692 15016 24704
rect 15068 24692 15074 24744
rect 15764 24704 17356 24732
rect 13262 24664 13268 24676
rect 13223 24636 13268 24664
rect 13262 24624 13268 24636
rect 13320 24624 13326 24676
rect 14274 24624 14280 24676
rect 14332 24664 14338 24676
rect 14461 24667 14519 24673
rect 14461 24664 14473 24667
rect 14332 24636 14473 24664
rect 14332 24624 14338 24636
rect 14461 24633 14473 24636
rect 14507 24633 14519 24667
rect 15764 24664 15792 24704
rect 17218 24664 17224 24676
rect 14461 24627 14519 24633
rect 15580 24636 15792 24664
rect 17179 24636 17224 24664
rect 12805 24599 12863 24605
rect 12805 24565 12817 24599
rect 12851 24596 12863 24599
rect 15580 24596 15608 24636
rect 17218 24624 17224 24636
rect 17276 24624 17282 24676
rect 17328 24664 17356 24704
rect 17494 24692 17500 24744
rect 17552 24732 17558 24744
rect 17681 24735 17739 24741
rect 17681 24732 17693 24735
rect 17552 24704 17693 24732
rect 17552 24692 17558 24704
rect 17681 24701 17693 24704
rect 17727 24701 17739 24735
rect 17681 24695 17739 24701
rect 17865 24735 17923 24741
rect 17865 24701 17877 24735
rect 17911 24732 17923 24735
rect 17954 24732 17960 24744
rect 17911 24704 17960 24732
rect 17911 24701 17923 24704
rect 17865 24695 17923 24701
rect 17954 24692 17960 24704
rect 18012 24692 18018 24744
rect 18509 24735 18567 24741
rect 18509 24701 18521 24735
rect 18555 24732 18567 24735
rect 19245 24735 19303 24741
rect 19245 24732 19257 24735
rect 18555 24704 19257 24732
rect 18555 24701 18567 24704
rect 18509 24695 18567 24701
rect 19245 24701 19257 24704
rect 19291 24732 19303 24735
rect 19610 24732 19616 24744
rect 19291 24704 19616 24732
rect 19291 24701 19303 24704
rect 19245 24695 19303 24701
rect 19610 24692 19616 24704
rect 19668 24732 19674 24744
rect 20070 24732 20076 24744
rect 19668 24704 20076 24732
rect 19668 24692 19674 24704
rect 20070 24692 20076 24704
rect 20128 24692 20134 24744
rect 20162 24692 20168 24744
rect 20220 24732 20226 24744
rect 20349 24735 20407 24741
rect 20220 24704 20265 24732
rect 20220 24692 20226 24704
rect 20349 24701 20361 24735
rect 20395 24732 20407 24735
rect 20622 24732 20628 24744
rect 20395 24704 20628 24732
rect 20395 24701 20407 24704
rect 20349 24695 20407 24701
rect 20622 24692 20628 24704
rect 20680 24732 20686 24744
rect 21266 24732 21272 24744
rect 20680 24704 21272 24732
rect 20680 24692 20686 24704
rect 21266 24692 21272 24704
rect 21324 24692 21330 24744
rect 23474 24692 23480 24744
rect 23532 24732 23538 24744
rect 24305 24735 24363 24741
rect 24305 24732 24317 24735
rect 23532 24704 24317 24732
rect 23532 24692 23538 24704
rect 24305 24701 24317 24704
rect 24351 24701 24363 24735
rect 24305 24695 24363 24701
rect 17328 24636 19288 24664
rect 12851 24568 15608 24596
rect 19260 24596 19288 24636
rect 20714 24624 20720 24676
rect 20772 24664 20778 24676
rect 20809 24667 20867 24673
rect 20809 24664 20821 24667
rect 20772 24636 20821 24664
rect 20772 24624 20778 24636
rect 20809 24633 20821 24636
rect 20855 24633 20867 24667
rect 20809 24627 20867 24633
rect 21174 24624 21180 24676
rect 21232 24664 21238 24676
rect 25424 24664 25452 24772
rect 28822 24769 28834 24772
rect 28868 24769 28880 24803
rect 28822 24763 28880 24769
rect 29089 24803 29147 24809
rect 29089 24769 29101 24803
rect 29135 24800 29147 24803
rect 29270 24800 29276 24812
rect 29135 24772 29276 24800
rect 29135 24769 29147 24772
rect 29089 24763 29147 24769
rect 29270 24760 29276 24772
rect 29328 24760 29334 24812
rect 29546 24800 29552 24812
rect 29507 24772 29552 24800
rect 29546 24760 29552 24772
rect 29604 24760 29610 24812
rect 31202 24800 31208 24812
rect 31163 24772 31208 24800
rect 31202 24760 31208 24772
rect 31260 24760 31266 24812
rect 32122 24760 32128 24812
rect 32180 24800 32186 24812
rect 33045 24803 33103 24809
rect 33045 24800 33057 24803
rect 32180 24772 33057 24800
rect 32180 24760 32186 24772
rect 33045 24769 33057 24772
rect 33091 24769 33103 24803
rect 33045 24763 33103 24769
rect 33134 24760 33140 24812
rect 33192 24800 33198 24812
rect 35161 24803 35219 24809
rect 35161 24800 35173 24803
rect 33192 24772 35173 24800
rect 33192 24760 33198 24772
rect 35161 24769 35173 24772
rect 35207 24769 35219 24803
rect 35161 24763 35219 24769
rect 35342 24760 35348 24812
rect 35400 24800 35406 24812
rect 35989 24803 36047 24809
rect 35989 24800 36001 24803
rect 35400 24772 36001 24800
rect 35400 24760 35406 24772
rect 35989 24769 36001 24772
rect 36035 24769 36047 24803
rect 37645 24803 37703 24809
rect 37645 24800 37657 24803
rect 35989 24763 36047 24769
rect 36740 24772 37657 24800
rect 29178 24692 29184 24744
rect 29236 24732 29242 24744
rect 34514 24732 34520 24744
rect 29236 24704 34520 24732
rect 29236 24692 29242 24704
rect 34514 24692 34520 24704
rect 34572 24692 34578 24744
rect 36740 24732 36768 24772
rect 37645 24769 37657 24772
rect 37691 24769 37703 24803
rect 37645 24763 37703 24769
rect 34624 24704 36768 24732
rect 27706 24664 27712 24676
rect 21232 24636 25452 24664
rect 27667 24636 27712 24664
rect 21232 24624 21238 24636
rect 27706 24624 27712 24636
rect 27764 24624 27770 24676
rect 29730 24664 29736 24676
rect 29691 24636 29736 24664
rect 29730 24624 29736 24636
rect 29788 24624 29794 24676
rect 31386 24664 31392 24676
rect 31347 24636 31392 24664
rect 31386 24624 31392 24636
rect 31444 24624 31450 24676
rect 33226 24664 33232 24676
rect 33187 24636 33232 24664
rect 33226 24624 33232 24636
rect 33284 24624 33290 24676
rect 33778 24624 33784 24676
rect 33836 24664 33842 24676
rect 34624 24664 34652 24704
rect 36814 24692 36820 24744
rect 36872 24732 36878 24744
rect 37461 24735 37519 24741
rect 37461 24732 37473 24735
rect 36872 24704 37473 24732
rect 36872 24692 36878 24704
rect 37461 24701 37473 24704
rect 37507 24701 37519 24735
rect 37461 24695 37519 24701
rect 33836 24636 34652 24664
rect 35345 24667 35403 24673
rect 33836 24624 33842 24636
rect 35345 24633 35357 24667
rect 35391 24664 35403 24667
rect 35986 24664 35992 24676
rect 35391 24636 35992 24664
rect 35391 24633 35403 24636
rect 35345 24627 35403 24633
rect 35986 24624 35992 24636
rect 36044 24624 36050 24676
rect 36170 24664 36176 24676
rect 36131 24636 36176 24664
rect 36170 24624 36176 24636
rect 36228 24624 36234 24676
rect 37826 24664 37832 24676
rect 36556 24636 37832 24664
rect 23198 24596 23204 24608
rect 19260 24568 23204 24596
rect 12851 24565 12863 24568
rect 12805 24559 12863 24565
rect 23198 24556 23204 24568
rect 23256 24556 23262 24608
rect 23293 24599 23351 24605
rect 23293 24565 23305 24599
rect 23339 24596 23351 24599
rect 23382 24596 23388 24608
rect 23339 24568 23388 24596
rect 23339 24565 23351 24568
rect 23293 24559 23351 24565
rect 23382 24556 23388 24568
rect 23440 24556 23446 24608
rect 23566 24556 23572 24608
rect 23624 24596 23630 24608
rect 23753 24599 23811 24605
rect 23753 24596 23765 24599
rect 23624 24568 23765 24596
rect 23624 24556 23630 24568
rect 23753 24565 23765 24568
rect 23799 24565 23811 24599
rect 23753 24559 23811 24565
rect 29822 24556 29828 24608
rect 29880 24596 29886 24608
rect 30193 24599 30251 24605
rect 30193 24596 30205 24599
rect 29880 24568 30205 24596
rect 29880 24556 29886 24568
rect 30193 24565 30205 24568
rect 30239 24596 30251 24599
rect 31570 24596 31576 24608
rect 30239 24568 31576 24596
rect 30239 24565 30251 24568
rect 30193 24559 30251 24565
rect 31570 24556 31576 24568
rect 31628 24596 31634 24608
rect 32125 24599 32183 24605
rect 32125 24596 32137 24599
rect 31628 24568 32137 24596
rect 31628 24556 31634 24568
rect 32125 24565 32137 24568
rect 32171 24565 32183 24599
rect 32125 24559 32183 24565
rect 33594 24556 33600 24608
rect 33652 24596 33658 24608
rect 33689 24599 33747 24605
rect 33689 24596 33701 24599
rect 33652 24568 33701 24596
rect 33652 24556 33658 24568
rect 33689 24565 33701 24568
rect 33735 24565 33747 24599
rect 34330 24596 34336 24608
rect 34243 24568 34336 24596
rect 33689 24559 33747 24565
rect 34330 24556 34336 24568
rect 34388 24596 34394 24608
rect 36556 24596 36584 24636
rect 37826 24624 37832 24636
rect 37884 24624 37890 24676
rect 34388 24568 36584 24596
rect 36725 24599 36783 24605
rect 34388 24556 34394 24568
rect 36725 24565 36737 24599
rect 36771 24596 36783 24599
rect 36814 24596 36820 24608
rect 36771 24568 36820 24596
rect 36771 24565 36783 24568
rect 36725 24559 36783 24565
rect 36814 24556 36820 24568
rect 36872 24556 36878 24608
rect 37918 24556 37924 24608
rect 37976 24596 37982 24608
rect 38105 24599 38163 24605
rect 38105 24596 38117 24599
rect 37976 24568 38117 24596
rect 37976 24556 37982 24568
rect 38105 24565 38117 24568
rect 38151 24565 38163 24599
rect 38105 24559 38163 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 13630 24352 13636 24404
rect 13688 24392 13694 24404
rect 14277 24395 14335 24401
rect 14277 24392 14289 24395
rect 13688 24364 14289 24392
rect 13688 24352 13694 24364
rect 14277 24361 14289 24364
rect 14323 24361 14335 24395
rect 14277 24355 14335 24361
rect 17678 24352 17684 24404
rect 17736 24392 17742 24404
rect 17773 24395 17831 24401
rect 17773 24392 17785 24395
rect 17736 24364 17785 24392
rect 17736 24352 17742 24364
rect 17773 24361 17785 24364
rect 17819 24361 17831 24395
rect 21174 24392 21180 24404
rect 21135 24364 21180 24392
rect 17773 24355 17831 24361
rect 21174 24352 21180 24364
rect 21232 24352 21238 24404
rect 22094 24352 22100 24404
rect 22152 24392 22158 24404
rect 22152 24364 22197 24392
rect 22152 24352 22158 24364
rect 23382 24352 23388 24404
rect 23440 24392 23446 24404
rect 26418 24392 26424 24404
rect 23440 24364 26424 24392
rect 23440 24352 23446 24364
rect 26418 24352 26424 24364
rect 26476 24352 26482 24404
rect 28077 24395 28135 24401
rect 28077 24361 28089 24395
rect 28123 24392 28135 24395
rect 29178 24392 29184 24404
rect 28123 24364 29184 24392
rect 28123 24361 28135 24364
rect 28077 24355 28135 24361
rect 29178 24352 29184 24364
rect 29236 24352 29242 24404
rect 29546 24392 29552 24404
rect 29507 24364 29552 24392
rect 29546 24352 29552 24364
rect 29604 24352 29610 24404
rect 32122 24392 32128 24404
rect 32083 24364 32128 24392
rect 32122 24352 32128 24364
rect 32180 24352 32186 24404
rect 35434 24352 35440 24404
rect 35492 24392 35498 24404
rect 35529 24395 35587 24401
rect 35529 24392 35541 24395
rect 35492 24364 35541 24392
rect 35492 24352 35498 24364
rect 35529 24361 35541 24364
rect 35575 24361 35587 24395
rect 36538 24392 36544 24404
rect 36499 24364 36544 24392
rect 35529 24355 35587 24361
rect 36538 24352 36544 24364
rect 36596 24352 36602 24404
rect 38010 24352 38016 24404
rect 38068 24392 38074 24404
rect 38105 24395 38163 24401
rect 38105 24392 38117 24395
rect 38068 24364 38117 24392
rect 38068 24352 38074 24364
rect 38105 24361 38117 24364
rect 38151 24361 38163 24395
rect 38105 24355 38163 24361
rect 16114 24284 16120 24336
rect 16172 24324 16178 24336
rect 20070 24324 20076 24336
rect 16172 24296 20076 24324
rect 16172 24284 16178 24296
rect 20070 24284 20076 24296
rect 20128 24324 20134 24336
rect 20441 24327 20499 24333
rect 20441 24324 20453 24327
rect 20128 24296 20453 24324
rect 20128 24284 20134 24296
rect 20441 24293 20453 24296
rect 20487 24293 20499 24327
rect 24854 24324 24860 24336
rect 20441 24287 20499 24293
rect 22066 24296 24860 24324
rect 18325 24259 18383 24265
rect 18325 24225 18337 24259
rect 18371 24256 18383 24259
rect 19610 24256 19616 24268
rect 18371 24228 19616 24256
rect 18371 24225 18383 24228
rect 18325 24219 18383 24225
rect 19610 24216 19616 24228
rect 19668 24256 19674 24268
rect 22066 24256 22094 24296
rect 24854 24284 24860 24296
rect 24912 24284 24918 24336
rect 25038 24324 25044 24336
rect 24999 24296 25044 24324
rect 25038 24284 25044 24296
rect 25096 24284 25102 24336
rect 28813 24327 28871 24333
rect 28813 24293 28825 24327
rect 28859 24293 28871 24327
rect 28813 24287 28871 24293
rect 30561 24327 30619 24333
rect 30561 24293 30573 24327
rect 30607 24324 30619 24327
rect 32214 24324 32220 24336
rect 30607 24296 32220 24324
rect 30607 24293 30619 24296
rect 30561 24287 30619 24293
rect 19668 24228 22094 24256
rect 22741 24259 22799 24265
rect 19668 24216 19674 24228
rect 22741 24225 22753 24259
rect 22787 24256 22799 24259
rect 22830 24256 22836 24268
rect 22787 24228 22836 24256
rect 22787 24225 22799 24228
rect 22741 24219 22799 24225
rect 22830 24216 22836 24228
rect 22888 24256 22894 24268
rect 23382 24256 23388 24268
rect 22888 24228 23388 24256
rect 22888 24216 22894 24228
rect 23382 24216 23388 24228
rect 23440 24216 23446 24268
rect 26326 24256 26332 24268
rect 23676 24228 26332 24256
rect 18506 24188 18512 24200
rect 18467 24160 18512 24188
rect 18506 24148 18512 24160
rect 18564 24148 18570 24200
rect 19797 24191 19855 24197
rect 19797 24157 19809 24191
rect 19843 24188 19855 24191
rect 19886 24188 19892 24200
rect 19843 24160 19892 24188
rect 19843 24157 19855 24160
rect 19797 24151 19855 24157
rect 19886 24148 19892 24160
rect 19944 24148 19950 24200
rect 19981 24191 20039 24197
rect 19981 24157 19993 24191
rect 20027 24188 20039 24191
rect 20993 24191 21051 24197
rect 20993 24188 21005 24191
rect 20027 24160 21005 24188
rect 20027 24157 20039 24160
rect 19981 24151 20039 24157
rect 20993 24157 21005 24160
rect 21039 24157 21051 24191
rect 23676 24188 23704 24228
rect 26326 24216 26332 24228
rect 26384 24216 26390 24268
rect 28828 24256 28856 24287
rect 32214 24284 32220 24296
rect 32272 24284 32278 24336
rect 35710 24324 35716 24336
rect 34716 24296 35716 24324
rect 33226 24256 33232 24268
rect 28828 24228 33232 24256
rect 33226 24216 33232 24228
rect 33284 24216 33290 24268
rect 33413 24259 33471 24265
rect 33413 24225 33425 24259
rect 33459 24256 33471 24259
rect 34146 24256 34152 24268
rect 33459 24228 34152 24256
rect 33459 24225 33471 24228
rect 33413 24219 33471 24225
rect 34146 24216 34152 24228
rect 34204 24216 34210 24268
rect 20993 24151 21051 24157
rect 21100 24160 23704 24188
rect 18874 24080 18880 24132
rect 18932 24120 18938 24132
rect 21100 24120 21128 24160
rect 23750 24148 23756 24200
rect 23808 24188 23814 24200
rect 27893 24191 27951 24197
rect 27893 24188 27905 24191
rect 23808 24160 27905 24188
rect 23808 24148 23814 24160
rect 27893 24157 27905 24160
rect 27939 24157 27951 24191
rect 27893 24151 27951 24157
rect 28074 24148 28080 24200
rect 28132 24188 28138 24200
rect 28629 24191 28687 24197
rect 28629 24188 28641 24191
rect 28132 24160 28641 24188
rect 28132 24148 28138 24160
rect 28629 24157 28641 24160
rect 28675 24157 28687 24191
rect 28629 24151 28687 24157
rect 28902 24148 28908 24200
rect 28960 24188 28966 24200
rect 29733 24191 29791 24197
rect 29733 24188 29745 24191
rect 28960 24160 29745 24188
rect 28960 24148 28966 24160
rect 29733 24157 29745 24160
rect 29779 24157 29791 24191
rect 29733 24151 29791 24157
rect 29822 24148 29828 24200
rect 29880 24188 29886 24200
rect 29880 24160 29925 24188
rect 29880 24148 29886 24160
rect 30006 24148 30012 24200
rect 30064 24188 30070 24200
rect 30377 24191 30435 24197
rect 30377 24188 30389 24191
rect 30064 24160 30389 24188
rect 30064 24148 30070 24160
rect 30377 24157 30389 24160
rect 30423 24157 30435 24191
rect 31018 24188 31024 24200
rect 30979 24160 31024 24188
rect 30377 24151 30435 24157
rect 31018 24148 31024 24160
rect 31076 24148 31082 24200
rect 31570 24148 31576 24200
rect 31628 24188 31634 24200
rect 31757 24191 31815 24197
rect 31757 24188 31769 24191
rect 31628 24160 31769 24188
rect 31628 24148 31634 24160
rect 31757 24157 31769 24160
rect 31803 24157 31815 24191
rect 31757 24151 31815 24157
rect 31941 24191 31999 24197
rect 31941 24157 31953 24191
rect 31987 24188 31999 24191
rect 32030 24188 32036 24200
rect 31987 24160 32036 24188
rect 31987 24157 31999 24160
rect 31941 24151 31999 24157
rect 32030 24148 32036 24160
rect 32088 24148 32094 24200
rect 33137 24191 33195 24197
rect 33137 24157 33149 24191
rect 33183 24188 33195 24191
rect 34330 24188 34336 24200
rect 33183 24160 34336 24188
rect 33183 24157 33195 24160
rect 33137 24151 33195 24157
rect 34330 24148 34336 24160
rect 34388 24148 34394 24200
rect 34514 24148 34520 24200
rect 34572 24188 34578 24200
rect 34716 24197 34744 24296
rect 35710 24284 35716 24296
rect 35768 24324 35774 24336
rect 37001 24327 37059 24333
rect 37001 24324 37013 24327
rect 35768 24296 37013 24324
rect 35768 24284 35774 24296
rect 37001 24293 37013 24296
rect 37047 24293 37059 24327
rect 37001 24287 37059 24293
rect 34701 24191 34759 24197
rect 34701 24188 34713 24191
rect 34572 24160 34713 24188
rect 34572 24148 34578 24160
rect 34701 24157 34713 24160
rect 34747 24157 34759 24191
rect 34701 24151 34759 24157
rect 34790 24148 34796 24200
rect 34848 24188 34854 24200
rect 34885 24191 34943 24197
rect 34885 24188 34897 24191
rect 34848 24160 34897 24188
rect 34848 24148 34854 24160
rect 34885 24157 34897 24160
rect 34931 24157 34943 24191
rect 35710 24188 35716 24200
rect 35671 24160 35716 24188
rect 34885 24151 34943 24157
rect 35710 24148 35716 24160
rect 35768 24148 35774 24200
rect 36357 24191 36415 24197
rect 36357 24188 36369 24191
rect 35866 24160 36369 24188
rect 18932 24092 21128 24120
rect 18932 24080 18938 24092
rect 21818 24080 21824 24132
rect 21876 24120 21882 24132
rect 22557 24123 22615 24129
rect 22557 24120 22569 24123
rect 21876 24092 22569 24120
rect 21876 24080 21882 24092
rect 22557 24089 22569 24092
rect 22603 24089 22615 24123
rect 23658 24120 23664 24132
rect 22557 24083 22615 24089
rect 23216 24092 23664 24120
rect 9122 24012 9128 24064
rect 9180 24052 9186 24064
rect 11974 24052 11980 24064
rect 9180 24024 11980 24052
rect 9180 24012 9186 24024
rect 11974 24012 11980 24024
rect 12032 24052 12038 24064
rect 12529 24055 12587 24061
rect 12529 24052 12541 24055
rect 12032 24024 12541 24052
rect 12032 24012 12038 24024
rect 12529 24021 12541 24024
rect 12575 24021 12587 24055
rect 15286 24052 15292 24064
rect 15247 24024 15292 24052
rect 12529 24015 12587 24021
rect 15286 24012 15292 24024
rect 15344 24012 15350 24064
rect 17313 24055 17371 24061
rect 17313 24021 17325 24055
rect 17359 24052 17371 24055
rect 17494 24052 17500 24064
rect 17359 24024 17500 24052
rect 17359 24021 17371 24024
rect 17313 24015 17371 24021
rect 17494 24012 17500 24024
rect 17552 24012 17558 24064
rect 18690 24052 18696 24064
rect 18651 24024 18696 24052
rect 18690 24012 18696 24024
rect 18748 24012 18754 24064
rect 22465 24055 22523 24061
rect 22465 24021 22477 24055
rect 22511 24052 22523 24055
rect 23216 24052 23244 24092
rect 23658 24080 23664 24092
rect 23716 24080 23722 24132
rect 24854 24080 24860 24132
rect 24912 24120 24918 24132
rect 30834 24120 30840 24132
rect 24912 24092 30840 24120
rect 24912 24080 24918 24092
rect 30834 24080 30840 24092
rect 30892 24080 30898 24132
rect 34606 24120 34612 24132
rect 31726 24092 34612 24120
rect 22511 24024 23244 24052
rect 22511 24021 22523 24024
rect 22465 24015 22523 24021
rect 23382 24012 23388 24064
rect 23440 24052 23446 24064
rect 24489 24055 24547 24061
rect 24489 24052 24501 24055
rect 23440 24024 24501 24052
rect 23440 24012 23446 24024
rect 24489 24021 24501 24024
rect 24535 24052 24547 24055
rect 25498 24052 25504 24064
rect 24535 24024 25504 24052
rect 24535 24021 24547 24024
rect 24489 24015 24547 24021
rect 25498 24012 25504 24024
rect 25556 24052 25562 24064
rect 25593 24055 25651 24061
rect 25593 24052 25605 24055
rect 25556 24024 25605 24052
rect 25556 24012 25562 24024
rect 25593 24021 25605 24024
rect 25639 24052 25651 24055
rect 26142 24052 26148 24064
rect 25639 24024 26148 24052
rect 25639 24021 25651 24024
rect 25593 24015 25651 24021
rect 26142 24012 26148 24024
rect 26200 24012 26206 24064
rect 31205 24055 31263 24061
rect 31205 24021 31217 24055
rect 31251 24052 31263 24055
rect 31726 24052 31754 24092
rect 34606 24080 34612 24092
rect 34664 24080 34670 24132
rect 35069 24123 35127 24129
rect 35069 24089 35081 24123
rect 35115 24120 35127 24123
rect 35866 24120 35894 24160
rect 36357 24157 36369 24160
rect 36403 24157 36415 24191
rect 36357 24151 36415 24157
rect 36446 24148 36452 24200
rect 36504 24188 36510 24200
rect 37737 24191 37795 24197
rect 37737 24188 37749 24191
rect 36504 24160 37749 24188
rect 36504 24148 36510 24160
rect 37737 24157 37749 24160
rect 37783 24157 37795 24191
rect 37918 24188 37924 24200
rect 37879 24160 37924 24188
rect 37737 24151 37795 24157
rect 37918 24148 37924 24160
rect 37976 24148 37982 24200
rect 35115 24092 35894 24120
rect 35115 24089 35127 24092
rect 35069 24083 35127 24089
rect 31251 24024 31754 24052
rect 31251 24021 31263 24024
rect 31205 24015 31263 24021
rect 32674 24012 32680 24064
rect 32732 24052 32738 24064
rect 32769 24055 32827 24061
rect 32769 24052 32781 24055
rect 32732 24024 32781 24052
rect 32732 24012 32738 24024
rect 32769 24021 32781 24024
rect 32815 24021 32827 24055
rect 32769 24015 32827 24021
rect 33229 24055 33287 24061
rect 33229 24021 33241 24055
rect 33275 24052 33287 24055
rect 33594 24052 33600 24064
rect 33275 24024 33600 24052
rect 33275 24021 33287 24024
rect 33229 24015 33287 24021
rect 33594 24012 33600 24024
rect 33652 24012 33658 24064
rect 34057 24055 34115 24061
rect 34057 24021 34069 24055
rect 34103 24052 34115 24055
rect 34146 24052 34152 24064
rect 34103 24024 34152 24052
rect 34103 24021 34115 24024
rect 34057 24015 34115 24021
rect 34146 24012 34152 24024
rect 34204 24012 34210 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 17405 23851 17463 23857
rect 17405 23817 17417 23851
rect 17451 23848 17463 23851
rect 17586 23848 17592 23860
rect 17451 23820 17592 23848
rect 17451 23817 17463 23820
rect 17405 23811 17463 23817
rect 17586 23808 17592 23820
rect 17644 23808 17650 23860
rect 18874 23848 18880 23860
rect 18835 23820 18880 23848
rect 18874 23808 18880 23820
rect 18932 23808 18938 23860
rect 19334 23808 19340 23860
rect 19392 23848 19398 23860
rect 19613 23851 19671 23857
rect 19613 23848 19625 23851
rect 19392 23820 19625 23848
rect 19392 23808 19398 23820
rect 19613 23817 19625 23820
rect 19659 23817 19671 23851
rect 19613 23811 19671 23817
rect 19981 23851 20039 23857
rect 19981 23817 19993 23851
rect 20027 23848 20039 23851
rect 20070 23848 20076 23860
rect 20027 23820 20076 23848
rect 20027 23817 20039 23820
rect 19981 23811 20039 23817
rect 20070 23808 20076 23820
rect 20128 23808 20134 23860
rect 22189 23851 22247 23857
rect 22189 23817 22201 23851
rect 22235 23848 22247 23851
rect 22370 23848 22376 23860
rect 22235 23820 22376 23848
rect 22235 23817 22247 23820
rect 22189 23811 22247 23817
rect 22370 23808 22376 23820
rect 22428 23808 22434 23860
rect 22649 23851 22707 23857
rect 22649 23817 22661 23851
rect 22695 23848 22707 23851
rect 23566 23848 23572 23860
rect 22695 23820 23572 23848
rect 22695 23817 22707 23820
rect 22649 23811 22707 23817
rect 23566 23808 23572 23820
rect 23624 23808 23630 23860
rect 23750 23848 23756 23860
rect 23711 23820 23756 23848
rect 23750 23808 23756 23820
rect 23808 23808 23814 23860
rect 24765 23851 24823 23857
rect 24765 23817 24777 23851
rect 24811 23848 24823 23851
rect 28350 23848 28356 23860
rect 24811 23820 28356 23848
rect 24811 23817 24823 23820
rect 24765 23811 24823 23817
rect 28350 23808 28356 23820
rect 28408 23808 28414 23860
rect 30009 23851 30067 23857
rect 30009 23817 30021 23851
rect 30055 23848 30067 23851
rect 31018 23848 31024 23860
rect 30055 23820 31024 23848
rect 30055 23817 30067 23820
rect 30009 23811 30067 23817
rect 31018 23808 31024 23820
rect 31076 23808 31082 23860
rect 31202 23848 31208 23860
rect 31163 23820 31208 23848
rect 31202 23808 31208 23820
rect 31260 23808 31266 23860
rect 32861 23851 32919 23857
rect 32861 23817 32873 23851
rect 32907 23848 32919 23851
rect 33134 23848 33140 23860
rect 32907 23820 33140 23848
rect 32907 23817 32919 23820
rect 32861 23811 32919 23817
rect 33134 23808 33140 23820
rect 33192 23808 33198 23860
rect 34790 23848 34796 23860
rect 34751 23820 34796 23848
rect 34790 23808 34796 23820
rect 34848 23808 34854 23860
rect 22557 23783 22615 23789
rect 22557 23780 22569 23783
rect 12406 23752 22569 23780
rect 11790 23468 11796 23520
rect 11848 23508 11854 23520
rect 12406 23508 12434 23752
rect 22557 23749 22569 23752
rect 22603 23780 22615 23783
rect 25038 23780 25044 23792
rect 22603 23752 25044 23780
rect 22603 23749 22615 23752
rect 22557 23743 22615 23749
rect 25038 23740 25044 23752
rect 25096 23740 25102 23792
rect 25958 23780 25964 23792
rect 25919 23752 25964 23780
rect 25958 23740 25964 23752
rect 26016 23780 26022 23792
rect 26602 23780 26608 23792
rect 26016 23752 26608 23780
rect 26016 23740 26022 23752
rect 26602 23740 26608 23752
rect 26660 23740 26666 23792
rect 28721 23783 28779 23789
rect 28721 23749 28733 23783
rect 28767 23780 28779 23783
rect 30190 23780 30196 23792
rect 28767 23752 30196 23780
rect 28767 23749 28779 23752
rect 28721 23743 28779 23749
rect 30190 23740 30196 23752
rect 30248 23740 30254 23792
rect 34425 23783 34483 23789
rect 34425 23749 34437 23783
rect 34471 23780 34483 23783
rect 37734 23780 37740 23792
rect 34471 23752 37740 23780
rect 34471 23749 34483 23752
rect 34425 23743 34483 23749
rect 37734 23740 37740 23752
rect 37792 23740 37798 23792
rect 17037 23715 17095 23721
rect 17037 23681 17049 23715
rect 17083 23712 17095 23715
rect 18690 23712 18696 23724
rect 17083 23684 18000 23712
rect 18651 23684 18696 23712
rect 17083 23681 17095 23684
rect 17037 23675 17095 23681
rect 16761 23647 16819 23653
rect 16761 23613 16773 23647
rect 16807 23613 16819 23647
rect 16942 23644 16948 23656
rect 16903 23616 16948 23644
rect 16761 23607 16819 23613
rect 16776 23576 16804 23607
rect 16942 23604 16948 23616
rect 17000 23604 17006 23656
rect 17972 23653 18000 23684
rect 18690 23672 18696 23684
rect 18748 23672 18754 23724
rect 20073 23715 20131 23721
rect 20073 23681 20085 23715
rect 20119 23712 20131 23715
rect 21450 23712 21456 23724
rect 20119 23684 21456 23712
rect 20119 23681 20131 23684
rect 20073 23675 20131 23681
rect 21450 23672 21456 23684
rect 21508 23672 21514 23724
rect 23474 23712 23480 23724
rect 23435 23684 23480 23712
rect 23474 23672 23480 23684
rect 23532 23672 23538 23724
rect 23569 23715 23627 23721
rect 23569 23681 23581 23715
rect 23615 23681 23627 23715
rect 24578 23712 24584 23724
rect 24539 23684 24584 23712
rect 23569 23675 23627 23681
rect 17957 23647 18015 23653
rect 17957 23613 17969 23647
rect 18003 23644 18015 23647
rect 18782 23644 18788 23656
rect 18003 23616 18788 23644
rect 18003 23613 18015 23616
rect 17957 23607 18015 23613
rect 18782 23604 18788 23616
rect 18840 23604 18846 23656
rect 20162 23604 20168 23656
rect 20220 23644 20226 23656
rect 20257 23647 20315 23653
rect 20257 23644 20269 23647
rect 20220 23616 20269 23644
rect 20220 23604 20226 23616
rect 20257 23613 20269 23616
rect 20303 23644 20315 23647
rect 20622 23644 20628 23656
rect 20303 23616 20628 23644
rect 20303 23613 20315 23616
rect 20257 23607 20315 23613
rect 20622 23604 20628 23616
rect 20680 23604 20686 23656
rect 22830 23644 22836 23656
rect 22791 23616 22836 23644
rect 22830 23604 22836 23616
rect 22888 23604 22894 23656
rect 23584 23644 23612 23675
rect 24578 23672 24584 23684
rect 24636 23672 24642 23724
rect 28813 23715 28871 23721
rect 28813 23681 28825 23715
rect 28859 23712 28871 23715
rect 29546 23712 29552 23724
rect 28859 23684 29552 23712
rect 28859 23681 28871 23684
rect 28813 23675 28871 23681
rect 29546 23672 29552 23684
rect 29604 23672 29610 23724
rect 29825 23715 29883 23721
rect 29825 23681 29837 23715
rect 29871 23712 29883 23715
rect 30650 23712 30656 23724
rect 29871 23684 30656 23712
rect 29871 23681 29883 23684
rect 29825 23675 29883 23681
rect 30650 23672 30656 23684
rect 30708 23672 30714 23724
rect 30834 23712 30840 23724
rect 30795 23684 30840 23712
rect 30834 23672 30840 23684
rect 30892 23672 30898 23724
rect 31018 23712 31024 23724
rect 30979 23684 31024 23712
rect 31018 23672 31024 23684
rect 31076 23672 31082 23724
rect 32674 23712 32680 23724
rect 32635 23684 32680 23712
rect 32674 23672 32680 23684
rect 32732 23672 32738 23724
rect 34514 23712 34520 23724
rect 33336 23684 34520 23712
rect 26050 23644 26056 23656
rect 23032 23616 23612 23644
rect 26011 23616 26056 23644
rect 20180 23576 20208 23604
rect 23032 23588 23060 23616
rect 26050 23604 26056 23616
rect 26108 23604 26114 23656
rect 26142 23604 26148 23656
rect 26200 23644 26206 23656
rect 27893 23647 27951 23653
rect 27893 23644 27905 23647
rect 26200 23616 27905 23644
rect 26200 23604 26206 23616
rect 27893 23613 27905 23616
rect 27939 23644 27951 23647
rect 28905 23647 28963 23653
rect 28905 23644 28917 23647
rect 27939 23616 28917 23644
rect 27939 23613 27951 23616
rect 27893 23607 27951 23613
rect 28905 23613 28917 23616
rect 28951 23613 28963 23647
rect 29638 23644 29644 23656
rect 29599 23616 29644 23644
rect 28905 23607 28963 23613
rect 29638 23604 29644 23616
rect 29696 23604 29702 23656
rect 30852 23644 30880 23672
rect 32490 23644 32496 23656
rect 30852 23616 32496 23644
rect 32490 23604 32496 23616
rect 32548 23644 32554 23656
rect 33336 23653 33364 23684
rect 34514 23672 34520 23684
rect 34572 23712 34578 23724
rect 35253 23715 35311 23721
rect 35253 23712 35265 23715
rect 34572 23684 35265 23712
rect 34572 23672 34578 23684
rect 35253 23681 35265 23684
rect 35299 23712 35311 23715
rect 35805 23715 35863 23721
rect 35805 23712 35817 23715
rect 35299 23684 35817 23712
rect 35299 23681 35311 23684
rect 35253 23675 35311 23681
rect 35805 23681 35817 23684
rect 35851 23681 35863 23715
rect 35805 23675 35863 23681
rect 33321 23647 33379 23653
rect 33321 23644 33333 23647
rect 32548 23616 33333 23644
rect 32548 23604 32554 23616
rect 33321 23613 33333 23616
rect 33367 23613 33379 23647
rect 34146 23644 34152 23656
rect 34107 23616 34152 23644
rect 33321 23607 33379 23613
rect 34146 23604 34152 23616
rect 34204 23604 34210 23656
rect 34333 23647 34391 23653
rect 34333 23613 34345 23647
rect 34379 23644 34391 23647
rect 34379 23616 35894 23644
rect 34379 23613 34391 23616
rect 34333 23607 34391 23613
rect 23014 23576 23020 23588
rect 16776 23548 20208 23576
rect 20272 23548 23020 23576
rect 11848 23480 12434 23508
rect 11848 23468 11854 23480
rect 19058 23468 19064 23520
rect 19116 23508 19122 23520
rect 20272 23508 20300 23548
rect 23014 23536 23020 23548
rect 23072 23536 23078 23588
rect 24670 23536 24676 23588
rect 24728 23576 24734 23588
rect 25593 23579 25651 23585
rect 25593 23576 25605 23579
rect 24728 23548 25605 23576
rect 24728 23536 24734 23548
rect 25593 23545 25605 23548
rect 25639 23545 25651 23579
rect 26068 23576 26096 23604
rect 26973 23579 27031 23585
rect 26973 23576 26985 23579
rect 26068 23548 26985 23576
rect 25593 23539 25651 23545
rect 26973 23545 26985 23548
rect 27019 23545 27031 23579
rect 26973 23539 27031 23545
rect 21174 23508 21180 23520
rect 19116 23480 20300 23508
rect 21135 23480 21180 23508
rect 19116 23468 19122 23480
rect 21174 23468 21180 23480
rect 21232 23468 21238 23520
rect 28258 23468 28264 23520
rect 28316 23508 28322 23520
rect 28353 23511 28411 23517
rect 28353 23508 28365 23511
rect 28316 23480 28365 23508
rect 28316 23468 28322 23480
rect 28353 23477 28365 23480
rect 28399 23477 28411 23511
rect 35866 23508 35894 23616
rect 36449 23511 36507 23517
rect 36449 23508 36461 23511
rect 35866 23480 36461 23508
rect 28353 23471 28411 23477
rect 36449 23477 36461 23480
rect 36495 23508 36507 23511
rect 37090 23508 37096 23520
rect 36495 23480 37096 23508
rect 36495 23477 36507 23480
rect 36449 23471 36507 23477
rect 37090 23468 37096 23480
rect 37148 23468 37154 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 16942 23264 16948 23316
rect 17000 23304 17006 23316
rect 17402 23304 17408 23316
rect 17000 23276 17408 23304
rect 17000 23264 17006 23276
rect 17402 23264 17408 23276
rect 17460 23304 17466 23316
rect 17497 23307 17555 23313
rect 17497 23304 17509 23307
rect 17460 23276 17509 23304
rect 17460 23264 17466 23276
rect 17497 23273 17509 23276
rect 17543 23273 17555 23307
rect 17497 23267 17555 23273
rect 21085 23307 21143 23313
rect 21085 23273 21097 23307
rect 21131 23304 21143 23307
rect 22002 23304 22008 23316
rect 21131 23276 22008 23304
rect 21131 23273 21143 23276
rect 21085 23267 21143 23273
rect 22002 23264 22008 23276
rect 22060 23264 22066 23316
rect 24578 23264 24584 23316
rect 24636 23304 24642 23316
rect 24765 23307 24823 23313
rect 24765 23304 24777 23307
rect 24636 23276 24777 23304
rect 24636 23264 24642 23276
rect 24765 23273 24777 23276
rect 24811 23273 24823 23307
rect 26602 23304 26608 23316
rect 26563 23276 26608 23304
rect 24765 23267 24823 23273
rect 26602 23264 26608 23276
rect 26660 23264 26666 23316
rect 29270 23264 29276 23316
rect 29328 23304 29334 23316
rect 29546 23304 29552 23316
rect 29328 23276 29552 23304
rect 29328 23264 29334 23276
rect 29546 23264 29552 23276
rect 29604 23264 29610 23316
rect 30190 23304 30196 23316
rect 30151 23276 30196 23304
rect 30190 23264 30196 23276
rect 30248 23264 30254 23316
rect 31754 23304 31760 23316
rect 31715 23276 31760 23304
rect 31754 23264 31760 23276
rect 31812 23264 31818 23316
rect 32490 23304 32496 23316
rect 32451 23276 32496 23304
rect 32490 23264 32496 23276
rect 32548 23264 32554 23316
rect 34698 23304 34704 23316
rect 34659 23276 34704 23304
rect 34698 23264 34704 23276
rect 34756 23264 34762 23316
rect 35529 23307 35587 23313
rect 35529 23273 35541 23307
rect 35575 23304 35587 23307
rect 35710 23304 35716 23316
rect 35575 23276 35716 23304
rect 35575 23273 35587 23276
rect 35529 23267 35587 23273
rect 35710 23264 35716 23276
rect 35768 23264 35774 23316
rect 35894 23264 35900 23316
rect 35952 23304 35958 23316
rect 36817 23307 36875 23313
rect 36817 23304 36829 23307
rect 35952 23276 36829 23304
rect 35952 23264 35958 23276
rect 36817 23273 36829 23276
rect 36863 23273 36875 23307
rect 36817 23267 36875 23273
rect 20346 23236 20352 23248
rect 19720 23208 20352 23236
rect 19720 23177 19748 23208
rect 20346 23196 20352 23208
rect 20404 23236 20410 23248
rect 33321 23239 33379 23245
rect 20404 23208 31754 23236
rect 20404 23196 20410 23208
rect 19705 23171 19763 23177
rect 19705 23137 19717 23171
rect 19751 23137 19763 23171
rect 19705 23131 19763 23137
rect 20533 23171 20591 23177
rect 20533 23137 20545 23171
rect 20579 23168 20591 23171
rect 20622 23168 20628 23180
rect 20579 23140 20628 23168
rect 20579 23137 20591 23140
rect 20533 23131 20591 23137
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23100 19947 23103
rect 20548 23100 20576 23131
rect 20622 23128 20628 23140
rect 20680 23128 20686 23180
rect 22281 23171 22339 23177
rect 22281 23168 22293 23171
rect 20732 23140 22293 23168
rect 20732 23109 20760 23140
rect 22281 23137 22293 23140
rect 22327 23168 22339 23171
rect 25866 23168 25872 23180
rect 22327 23140 25872 23168
rect 22327 23137 22339 23140
rect 22281 23131 22339 23137
rect 25866 23128 25872 23140
rect 25924 23128 25930 23180
rect 28997 23171 29055 23177
rect 28997 23168 29009 23171
rect 25976 23140 29009 23168
rect 19935 23072 20576 23100
rect 20717 23103 20775 23109
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 20717 23069 20729 23103
rect 20763 23069 20775 23103
rect 23014 23100 23020 23112
rect 22975 23072 23020 23100
rect 20717 23063 20775 23069
rect 23014 23060 23020 23072
rect 23072 23100 23078 23112
rect 23661 23103 23719 23109
rect 23661 23100 23673 23103
rect 23072 23072 23673 23100
rect 23072 23060 23078 23072
rect 23661 23069 23673 23072
rect 23707 23100 23719 23103
rect 23842 23100 23848 23112
rect 23707 23072 23848 23100
rect 23707 23069 23719 23072
rect 23661 23063 23719 23069
rect 23842 23060 23848 23072
rect 23900 23060 23906 23112
rect 24489 23103 24547 23109
rect 24489 23069 24501 23103
rect 24535 23069 24547 23103
rect 24489 23063 24547 23069
rect 24581 23103 24639 23109
rect 24581 23069 24593 23103
rect 24627 23100 24639 23103
rect 24670 23100 24676 23112
rect 24627 23072 24676 23100
rect 24627 23069 24639 23072
rect 24581 23063 24639 23069
rect 20625 23035 20683 23041
rect 20625 23001 20637 23035
rect 20671 23032 20683 23035
rect 20806 23032 20812 23044
rect 20671 23004 20812 23032
rect 20671 23001 20683 23004
rect 20625 22995 20683 23001
rect 20806 22992 20812 23004
rect 20864 23032 20870 23044
rect 21174 23032 21180 23044
rect 20864 23004 21180 23032
rect 20864 22992 20870 23004
rect 21174 22992 21180 23004
rect 21232 22992 21238 23044
rect 22830 23032 22836 23044
rect 22066 23004 22836 23032
rect 21726 22964 21732 22976
rect 21687 22936 21732 22964
rect 21726 22924 21732 22936
rect 21784 22964 21790 22976
rect 22066 22964 22094 23004
rect 22830 22992 22836 23004
rect 22888 22992 22894 23044
rect 24504 23032 24532 23063
rect 24670 23060 24676 23072
rect 24728 23060 24734 23112
rect 25222 23100 25228 23112
rect 25183 23072 25228 23100
rect 25222 23060 25228 23072
rect 25280 23060 25286 23112
rect 25976 23100 26004 23140
rect 28997 23137 29009 23140
rect 29043 23168 29055 23171
rect 29638 23168 29644 23180
rect 29043 23140 29644 23168
rect 29043 23137 29055 23140
rect 28997 23131 29055 23137
rect 29638 23128 29644 23140
rect 29696 23128 29702 23180
rect 31726 23168 31754 23208
rect 33321 23205 33333 23239
rect 33367 23236 33379 23239
rect 35342 23236 35348 23248
rect 33367 23208 35348 23236
rect 33367 23205 33379 23208
rect 33321 23199 33379 23205
rect 35342 23196 35348 23208
rect 35400 23196 35406 23248
rect 33873 23171 33931 23177
rect 33873 23168 33885 23171
rect 31726 23140 33885 23168
rect 33873 23137 33885 23140
rect 33919 23168 33931 23171
rect 34146 23168 34152 23180
rect 33919 23140 34152 23168
rect 33919 23137 33931 23140
rect 33873 23131 33931 23137
rect 34146 23128 34152 23140
rect 34204 23128 34210 23180
rect 34514 23128 34520 23180
rect 34572 23168 34578 23180
rect 35069 23171 35127 23177
rect 35069 23168 35081 23171
rect 34572 23140 35081 23168
rect 34572 23128 34578 23140
rect 35069 23137 35081 23140
rect 35115 23168 35127 23171
rect 35897 23171 35955 23177
rect 35897 23168 35909 23171
rect 35115 23140 35909 23168
rect 35115 23137 35127 23140
rect 35069 23131 35127 23137
rect 35897 23137 35909 23140
rect 35943 23137 35955 23171
rect 35897 23131 35955 23137
rect 28258 23100 28264 23112
rect 25332 23072 26004 23100
rect 28219 23072 28264 23100
rect 25332 23032 25360 23072
rect 28258 23060 28264 23072
rect 28316 23060 28322 23112
rect 28445 23103 28503 23109
rect 28445 23069 28457 23103
rect 28491 23100 28503 23103
rect 30374 23100 30380 23112
rect 28491 23072 30380 23100
rect 28491 23069 28503 23072
rect 28445 23063 28503 23069
rect 30374 23060 30380 23072
rect 30432 23100 30438 23112
rect 30745 23103 30803 23109
rect 30745 23100 30757 23103
rect 30432 23072 30757 23100
rect 30432 23060 30438 23072
rect 30745 23069 30757 23072
rect 30791 23069 30803 23103
rect 30926 23100 30932 23112
rect 30887 23072 30932 23100
rect 30745 23063 30803 23069
rect 30926 23060 30932 23072
rect 30984 23060 30990 23112
rect 31113 23103 31171 23109
rect 31113 23069 31125 23103
rect 31159 23100 31171 23103
rect 31573 23103 31631 23109
rect 31573 23100 31585 23103
rect 31159 23072 31585 23100
rect 31159 23069 31171 23072
rect 31113 23063 31171 23069
rect 31573 23069 31585 23072
rect 31619 23069 31631 23103
rect 31573 23063 31631 23069
rect 32490 23060 32496 23112
rect 32548 23100 32554 23112
rect 32953 23103 33011 23109
rect 32953 23100 32965 23103
rect 32548 23072 32965 23100
rect 32548 23060 32554 23072
rect 32953 23069 32965 23072
rect 32999 23069 33011 23103
rect 33134 23100 33140 23112
rect 33095 23072 33140 23100
rect 32953 23063 33011 23069
rect 33134 23060 33140 23072
rect 33192 23060 33198 23112
rect 34882 23100 34888 23112
rect 34843 23072 34888 23100
rect 34882 23060 34888 23072
rect 34940 23060 34946 23112
rect 35713 23103 35771 23109
rect 35713 23069 35725 23103
rect 35759 23100 35771 23103
rect 36998 23100 37004 23112
rect 35759 23072 35894 23100
rect 36959 23072 37004 23100
rect 35759 23069 35771 23072
rect 35713 23063 35771 23069
rect 31846 23032 31852 23044
rect 24504 23004 25360 23032
rect 25424 23004 31852 23032
rect 23106 22964 23112 22976
rect 21784 22936 22094 22964
rect 23067 22936 23112 22964
rect 21784 22924 21790 22936
rect 23106 22924 23112 22936
rect 23164 22924 23170 22976
rect 24394 22924 24400 22976
rect 24452 22964 24458 22976
rect 24504 22964 24532 23004
rect 25424 22973 25452 23004
rect 31846 22992 31852 23004
rect 31904 22992 31910 23044
rect 35866 22976 35894 23072
rect 36998 23060 37004 23072
rect 37056 23060 37062 23112
rect 24452 22936 24532 22964
rect 25409 22967 25467 22973
rect 24452 22924 24458 22936
rect 25409 22933 25421 22967
rect 25455 22933 25467 22967
rect 25409 22927 25467 22933
rect 27706 22924 27712 22976
rect 27764 22964 27770 22976
rect 28077 22967 28135 22973
rect 28077 22964 28089 22967
rect 27764 22936 28089 22964
rect 27764 22924 27770 22936
rect 28077 22933 28089 22936
rect 28123 22933 28135 22967
rect 35866 22936 35900 22976
rect 28077 22927 28135 22933
rect 35894 22924 35900 22936
rect 35952 22924 35958 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 23106 22720 23112 22772
rect 23164 22720 23170 22772
rect 23385 22763 23443 22769
rect 23385 22729 23397 22763
rect 23431 22760 23443 22763
rect 25222 22760 25228 22772
rect 23431 22732 25228 22760
rect 23431 22729 23443 22732
rect 23385 22723 23443 22729
rect 25222 22720 25228 22732
rect 25280 22720 25286 22772
rect 28537 22763 28595 22769
rect 28537 22729 28549 22763
rect 28583 22729 28595 22763
rect 30006 22760 30012 22772
rect 29967 22732 30012 22760
rect 28537 22723 28595 22729
rect 23124 22692 23152 22720
rect 23842 22692 23848 22704
rect 23032 22664 23336 22692
rect 23803 22664 23848 22692
rect 20622 22584 20628 22636
rect 20680 22624 20686 22636
rect 20809 22627 20867 22633
rect 20809 22624 20821 22627
rect 20680 22596 20821 22624
rect 20680 22584 20686 22596
rect 20809 22593 20821 22596
rect 20855 22624 20867 22627
rect 21818 22624 21824 22636
rect 20855 22596 21824 22624
rect 20855 22593 20867 22596
rect 20809 22587 20867 22593
rect 21818 22584 21824 22596
rect 21876 22584 21882 22636
rect 22189 22627 22247 22633
rect 22189 22593 22201 22627
rect 22235 22624 22247 22627
rect 22554 22624 22560 22636
rect 22235 22596 22560 22624
rect 22235 22593 22247 22596
rect 22189 22587 22247 22593
rect 22554 22584 22560 22596
rect 22612 22584 22618 22636
rect 23032 22633 23060 22664
rect 23017 22627 23075 22633
rect 23017 22593 23029 22627
rect 23063 22593 23075 22627
rect 23017 22587 23075 22593
rect 23201 22627 23259 22633
rect 23201 22593 23213 22627
rect 23247 22593 23259 22627
rect 23201 22587 23259 22593
rect 21085 22559 21143 22565
rect 21085 22525 21097 22559
rect 21131 22556 21143 22559
rect 21726 22556 21732 22568
rect 21131 22528 21732 22556
rect 21131 22525 21143 22528
rect 21085 22519 21143 22525
rect 21726 22516 21732 22528
rect 21784 22556 21790 22568
rect 21913 22559 21971 22565
rect 21913 22556 21925 22559
rect 21784 22528 21925 22556
rect 21784 22516 21790 22528
rect 21913 22525 21925 22528
rect 21959 22525 21971 22559
rect 21913 22519 21971 22525
rect 22094 22516 22100 22568
rect 22152 22556 22158 22568
rect 22152 22528 22197 22556
rect 22152 22516 22158 22528
rect 22557 22491 22615 22497
rect 22557 22457 22569 22491
rect 22603 22488 22615 22491
rect 23216 22488 23244 22587
rect 23308 22556 23336 22664
rect 23842 22652 23848 22664
rect 23900 22652 23906 22704
rect 24394 22692 24400 22704
rect 24355 22664 24400 22692
rect 24394 22652 24400 22664
rect 24452 22652 24458 22704
rect 28552 22692 28580 22723
rect 30006 22720 30012 22732
rect 30064 22720 30070 22772
rect 30745 22763 30803 22769
rect 30745 22729 30757 22763
rect 30791 22760 30803 22763
rect 30834 22760 30840 22772
rect 30791 22732 30840 22760
rect 30791 22729 30803 22732
rect 30745 22723 30803 22729
rect 30834 22720 30840 22732
rect 30892 22720 30898 22772
rect 32306 22760 32312 22772
rect 32267 22732 32312 22760
rect 32306 22720 32312 22732
rect 32364 22720 32370 22772
rect 32490 22720 32496 22772
rect 32548 22760 32554 22772
rect 33321 22763 33379 22769
rect 33321 22760 33333 22763
rect 32548 22732 33333 22760
rect 32548 22720 32554 22732
rect 33321 22729 33333 22732
rect 33367 22729 33379 22763
rect 33321 22723 33379 22729
rect 30558 22692 30564 22704
rect 28552 22664 30564 22692
rect 30558 22652 30564 22664
rect 30616 22652 30622 22704
rect 25590 22624 25596 22636
rect 25551 22596 25596 22624
rect 25590 22584 25596 22596
rect 25648 22584 25654 22636
rect 25777 22627 25835 22633
rect 25777 22593 25789 22627
rect 25823 22624 25835 22627
rect 27065 22627 27123 22633
rect 27065 22624 27077 22627
rect 25823 22596 27077 22624
rect 25823 22593 25835 22596
rect 25777 22587 25835 22593
rect 27065 22593 27077 22596
rect 27111 22593 27123 22627
rect 27706 22624 27712 22636
rect 27667 22596 27712 22624
rect 27065 22587 27123 22593
rect 27706 22584 27712 22596
rect 27764 22584 27770 22636
rect 28350 22624 28356 22636
rect 28311 22596 28356 22624
rect 28350 22584 28356 22596
rect 28408 22584 28414 22636
rect 29822 22624 29828 22636
rect 29783 22596 29828 22624
rect 29822 22584 29828 22596
rect 29880 22584 29886 22636
rect 30190 22584 30196 22636
rect 30248 22624 30254 22636
rect 32125 22627 32183 22633
rect 32125 22624 32137 22627
rect 30248 22596 32137 22624
rect 30248 22584 30254 22596
rect 32125 22593 32137 22596
rect 32171 22593 32183 22627
rect 32125 22587 32183 22593
rect 25409 22559 25467 22565
rect 25409 22556 25421 22559
rect 23308 22528 25421 22556
rect 25409 22525 25421 22528
rect 25455 22556 25467 22559
rect 27614 22556 27620 22568
rect 25455 22528 27620 22556
rect 25455 22525 25467 22528
rect 25409 22519 25467 22525
rect 27614 22516 27620 22528
rect 27672 22516 27678 22568
rect 29641 22559 29699 22565
rect 29641 22525 29653 22559
rect 29687 22556 29699 22559
rect 30374 22556 30380 22568
rect 29687 22528 30380 22556
rect 29687 22525 29699 22528
rect 29641 22519 29699 22525
rect 30374 22516 30380 22528
rect 30432 22516 30438 22568
rect 33336 22556 33364 22723
rect 33686 22720 33692 22772
rect 33744 22760 33750 22772
rect 33873 22763 33931 22769
rect 33873 22760 33885 22763
rect 33744 22732 33885 22760
rect 33744 22720 33750 22732
rect 33873 22729 33885 22732
rect 33919 22729 33931 22763
rect 33873 22723 33931 22729
rect 34882 22720 34888 22772
rect 34940 22760 34946 22772
rect 35253 22763 35311 22769
rect 35253 22760 35265 22763
rect 34940 22732 35265 22760
rect 34940 22720 34946 22732
rect 35253 22729 35265 22732
rect 35299 22729 35311 22763
rect 35253 22723 35311 22729
rect 35621 22763 35679 22769
rect 35621 22729 35633 22763
rect 35667 22760 35679 22763
rect 36354 22760 36360 22772
rect 35667 22732 36360 22760
rect 35667 22729 35679 22732
rect 35621 22723 35679 22729
rect 36354 22720 36360 22732
rect 36412 22720 36418 22772
rect 35710 22692 35716 22704
rect 35671 22664 35716 22692
rect 35710 22652 35716 22664
rect 35768 22652 35774 22704
rect 34057 22627 34115 22633
rect 34057 22593 34069 22627
rect 34103 22624 34115 22627
rect 34698 22624 34704 22636
rect 34103 22596 34704 22624
rect 34103 22593 34115 22596
rect 34057 22587 34115 22593
rect 34698 22584 34704 22596
rect 34756 22584 34762 22636
rect 34241 22559 34299 22565
rect 34241 22556 34253 22559
rect 33336 22528 34253 22556
rect 34241 22525 34253 22528
rect 34287 22525 34299 22559
rect 35802 22556 35808 22568
rect 35763 22528 35808 22556
rect 34241 22519 34299 22525
rect 35802 22516 35808 22528
rect 35860 22516 35866 22568
rect 22603 22460 23244 22488
rect 27893 22491 27951 22497
rect 22603 22457 22615 22460
rect 22557 22451 22615 22457
rect 27893 22457 27905 22491
rect 27939 22488 27951 22491
rect 30466 22488 30472 22500
rect 27939 22460 30472 22488
rect 27939 22457 27951 22460
rect 27893 22451 27951 22457
rect 30466 22448 30472 22460
rect 30524 22448 30530 22500
rect 30742 22488 30748 22500
rect 30576 22460 30748 22488
rect 27249 22423 27307 22429
rect 27249 22389 27261 22423
rect 27295 22420 27307 22423
rect 30576 22420 30604 22460
rect 30742 22448 30748 22460
rect 30800 22448 30806 22500
rect 27295 22392 30604 22420
rect 27295 22389 27307 22392
rect 27249 22383 27307 22389
rect 34606 22380 34612 22432
rect 34664 22420 34670 22432
rect 34701 22423 34759 22429
rect 34701 22420 34713 22423
rect 34664 22392 34713 22420
rect 34664 22380 34670 22392
rect 34701 22389 34713 22392
rect 34747 22420 34759 22423
rect 38102 22420 38108 22432
rect 34747 22392 38108 22420
rect 34747 22389 34759 22392
rect 34701 22383 34759 22389
rect 38102 22380 38108 22392
rect 38160 22380 38166 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 25590 22176 25596 22228
rect 25648 22216 25654 22228
rect 26145 22219 26203 22225
rect 26145 22216 26157 22219
rect 25648 22188 26157 22216
rect 25648 22176 25654 22188
rect 26145 22185 26157 22188
rect 26191 22185 26203 22219
rect 26145 22179 26203 22185
rect 28350 22176 28356 22228
rect 28408 22216 28414 22228
rect 28445 22219 28503 22225
rect 28445 22216 28457 22219
rect 28408 22188 28457 22216
rect 28408 22176 28414 22188
rect 28445 22185 28457 22188
rect 28491 22185 28503 22219
rect 28445 22179 28503 22185
rect 33134 22176 33140 22228
rect 33192 22216 33198 22228
rect 33413 22219 33471 22225
rect 33413 22216 33425 22219
rect 33192 22188 33425 22216
rect 33192 22176 33198 22188
rect 33413 22185 33425 22188
rect 33459 22185 33471 22219
rect 34698 22216 34704 22228
rect 34659 22188 34704 22216
rect 33413 22179 33471 22185
rect 34698 22176 34704 22188
rect 34756 22176 34762 22228
rect 35894 22176 35900 22228
rect 35952 22216 35958 22228
rect 35952 22188 35997 22216
rect 35952 22176 35958 22188
rect 10962 22108 10968 22160
rect 11020 22148 11026 22160
rect 11974 22148 11980 22160
rect 11020 22120 11980 22148
rect 11020 22108 11026 22120
rect 11974 22108 11980 22120
rect 12032 22108 12038 22160
rect 22554 22108 22560 22160
rect 22612 22148 22618 22160
rect 23293 22151 23351 22157
rect 23293 22148 23305 22151
rect 22612 22120 23305 22148
rect 22612 22108 22618 22120
rect 23293 22117 23305 22120
rect 23339 22148 23351 22151
rect 28166 22148 28172 22160
rect 23339 22120 28172 22148
rect 23339 22117 23351 22120
rect 23293 22111 23351 22117
rect 28166 22108 28172 22120
rect 28224 22108 28230 22160
rect 30374 22148 30380 22160
rect 29840 22120 30380 22148
rect 25498 22040 25504 22092
rect 25556 22080 25562 22092
rect 25593 22083 25651 22089
rect 25593 22080 25605 22083
rect 25556 22052 25605 22080
rect 25556 22040 25562 22052
rect 25593 22049 25605 22052
rect 25639 22080 25651 22083
rect 26786 22080 26792 22092
rect 25639 22052 26792 22080
rect 25639 22049 25651 22052
rect 25593 22043 25651 22049
rect 26786 22040 26792 22052
rect 26844 22040 26850 22092
rect 27614 22080 27620 22092
rect 27527 22052 27620 22080
rect 27614 22040 27620 22052
rect 27672 22080 27678 22092
rect 29840 22089 29868 22120
rect 30374 22108 30380 22120
rect 30432 22148 30438 22160
rect 31478 22148 31484 22160
rect 30432 22120 31484 22148
rect 30432 22108 30438 22120
rect 31478 22108 31484 22120
rect 31536 22108 31542 22160
rect 28813 22083 28871 22089
rect 28813 22080 28825 22083
rect 27672 22052 28825 22080
rect 27672 22040 27678 22052
rect 28813 22049 28825 22052
rect 28859 22080 28871 22083
rect 29825 22083 29883 22089
rect 29825 22080 29837 22083
rect 28859 22052 29837 22080
rect 28859 22049 28871 22052
rect 28813 22043 28871 22049
rect 29825 22049 29837 22052
rect 29871 22049 29883 22083
rect 30190 22080 30196 22092
rect 30151 22052 30196 22080
rect 29825 22043 29883 22049
rect 30190 22040 30196 22052
rect 30248 22040 30254 22092
rect 30282 22040 30288 22092
rect 30340 22080 30346 22092
rect 33965 22083 34023 22089
rect 33965 22080 33977 22083
rect 30340 22052 33977 22080
rect 30340 22040 30346 22052
rect 33965 22049 33977 22052
rect 34011 22080 34023 22083
rect 35253 22083 35311 22089
rect 35253 22080 35265 22083
rect 34011 22052 35265 22080
rect 34011 22049 34023 22052
rect 33965 22043 34023 22049
rect 35253 22049 35265 22052
rect 35299 22080 35311 22083
rect 35802 22080 35808 22092
rect 35299 22052 35808 22080
rect 35299 22049 35311 22052
rect 35253 22043 35311 22049
rect 35802 22040 35808 22052
rect 35860 22080 35866 22092
rect 36449 22083 36507 22089
rect 36449 22080 36461 22083
rect 35860 22052 36461 22080
rect 35860 22040 35866 22052
rect 36449 22049 36461 22052
rect 36495 22049 36507 22083
rect 36449 22043 36507 22049
rect 16390 21972 16396 22024
rect 16448 22012 16454 22024
rect 20346 22012 20352 22024
rect 16448 21984 20352 22012
rect 16448 21972 16454 21984
rect 20346 21972 20352 21984
rect 20404 21972 20410 22024
rect 21818 22012 21824 22024
rect 21779 21984 21824 22012
rect 21818 21972 21824 21984
rect 21876 21972 21882 22024
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22741 22015 22799 22021
rect 22741 22012 22753 22015
rect 22152 21984 22753 22012
rect 22152 21972 22158 21984
rect 22741 21981 22753 21984
rect 22787 22012 22799 22015
rect 26970 22012 26976 22024
rect 22787 21984 26976 22012
rect 22787 21981 22799 21984
rect 22741 21975 22799 21981
rect 26970 21972 26976 21984
rect 27028 21972 27034 22024
rect 27801 22015 27859 22021
rect 27801 21981 27813 22015
rect 27847 22012 27859 22015
rect 27982 22012 27988 22024
rect 27847 21984 27988 22012
rect 27847 21981 27859 21984
rect 27801 21975 27859 21981
rect 27982 21972 27988 21984
rect 28040 21972 28046 22024
rect 28626 22012 28632 22024
rect 28587 21984 28632 22012
rect 28626 21972 28632 21984
rect 28684 21972 28690 22024
rect 30006 22012 30012 22024
rect 29967 21984 30012 22012
rect 30006 21972 30012 21984
rect 30064 21972 30070 22024
rect 33781 22015 33839 22021
rect 33781 21981 33793 22015
rect 33827 22012 33839 22015
rect 34606 22012 34612 22024
rect 33827 21984 34612 22012
rect 33827 21981 33839 21984
rect 33781 21975 33839 21981
rect 34606 21972 34612 21984
rect 34664 21972 34670 22024
rect 35069 22015 35127 22021
rect 35069 21981 35081 22015
rect 35115 22012 35127 22015
rect 35618 22012 35624 22024
rect 35115 21984 35624 22012
rect 35115 21981 35127 21984
rect 35069 21975 35127 21981
rect 35618 21972 35624 21984
rect 35676 21972 35682 22024
rect 36262 22012 36268 22024
rect 36223 21984 36268 22012
rect 36262 21972 36268 21984
rect 36320 21972 36326 22024
rect 26513 21947 26571 21953
rect 26513 21913 26525 21947
rect 26559 21944 26571 21947
rect 27246 21944 27252 21956
rect 26559 21916 27252 21944
rect 26559 21913 26571 21916
rect 26513 21907 26571 21913
rect 27246 21904 27252 21916
rect 27304 21944 27310 21956
rect 30098 21944 30104 21956
rect 27304 21916 30104 21944
rect 27304 21904 27310 21916
rect 30098 21904 30104 21916
rect 30156 21904 30162 21956
rect 22094 21876 22100 21888
rect 22055 21848 22100 21876
rect 22094 21836 22100 21848
rect 22152 21836 22158 21888
rect 26605 21879 26663 21885
rect 26605 21845 26617 21879
rect 26651 21876 26663 21879
rect 27154 21876 27160 21888
rect 26651 21848 27160 21876
rect 26651 21845 26663 21848
rect 26605 21839 26663 21845
rect 27154 21836 27160 21848
rect 27212 21836 27218 21888
rect 27985 21879 28043 21885
rect 27985 21845 27997 21879
rect 28031 21876 28043 21879
rect 28074 21876 28080 21888
rect 28031 21848 28080 21876
rect 28031 21845 28043 21848
rect 27985 21839 28043 21845
rect 28074 21836 28080 21848
rect 28132 21836 28138 21888
rect 32766 21836 32772 21888
rect 32824 21876 32830 21888
rect 33873 21879 33931 21885
rect 33873 21876 33885 21879
rect 32824 21848 33885 21876
rect 32824 21836 32830 21848
rect 33873 21845 33885 21848
rect 33919 21845 33931 21879
rect 33873 21839 33931 21845
rect 35161 21879 35219 21885
rect 35161 21845 35173 21879
rect 35207 21876 35219 21879
rect 35434 21876 35440 21888
rect 35207 21848 35440 21876
rect 35207 21845 35219 21848
rect 35161 21839 35219 21845
rect 35434 21836 35440 21848
rect 35492 21836 35498 21888
rect 36357 21879 36415 21885
rect 36357 21845 36369 21879
rect 36403 21876 36415 21879
rect 37185 21879 37243 21885
rect 37185 21876 37197 21879
rect 36403 21848 37197 21876
rect 36403 21845 36415 21848
rect 36357 21839 36415 21845
rect 37185 21845 37197 21848
rect 37231 21876 37243 21879
rect 37366 21876 37372 21888
rect 37231 21848 37372 21876
rect 37231 21845 37243 21848
rect 37185 21839 37243 21845
rect 37366 21836 37372 21848
rect 37424 21836 37430 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 28626 21672 28632 21684
rect 28587 21644 28632 21672
rect 28626 21632 28632 21644
rect 28684 21632 28690 21684
rect 30837 21675 30895 21681
rect 30837 21641 30849 21675
rect 30883 21672 30895 21675
rect 31018 21672 31024 21684
rect 30883 21644 31024 21672
rect 30883 21641 30895 21644
rect 30837 21635 30895 21641
rect 31018 21632 31024 21644
rect 31076 21632 31082 21684
rect 31205 21675 31263 21681
rect 31205 21641 31217 21675
rect 31251 21672 31263 21675
rect 32769 21675 32827 21681
rect 32769 21672 32781 21675
rect 31251 21644 32781 21672
rect 31251 21641 31263 21644
rect 31205 21635 31263 21641
rect 32769 21641 32781 21644
rect 32815 21672 32827 21675
rect 34790 21672 34796 21684
rect 32815 21644 34796 21672
rect 32815 21641 32827 21644
rect 32769 21635 32827 21641
rect 34790 21632 34796 21644
rect 34848 21632 34854 21684
rect 36449 21675 36507 21681
rect 36449 21641 36461 21675
rect 36495 21672 36507 21675
rect 36998 21672 37004 21684
rect 36495 21644 37004 21672
rect 36495 21641 36507 21644
rect 36449 21635 36507 21641
rect 36998 21632 37004 21644
rect 37056 21632 37062 21684
rect 31297 21607 31355 21613
rect 31297 21573 31309 21607
rect 31343 21604 31355 21607
rect 31386 21604 31392 21616
rect 31343 21576 31392 21604
rect 31343 21573 31355 21576
rect 31297 21567 31355 21573
rect 31386 21564 31392 21576
rect 31444 21604 31450 21616
rect 32125 21607 32183 21613
rect 32125 21604 32137 21607
rect 31444 21576 32137 21604
rect 31444 21564 31450 21576
rect 32125 21573 32137 21576
rect 32171 21573 32183 21607
rect 32125 21567 32183 21573
rect 28261 21539 28319 21545
rect 28261 21505 28273 21539
rect 28307 21536 28319 21539
rect 30285 21539 30343 21545
rect 30285 21536 30297 21539
rect 28307 21508 30297 21536
rect 28307 21505 28319 21508
rect 28261 21499 28319 21505
rect 30285 21505 30297 21508
rect 30331 21536 30343 21539
rect 32858 21536 32864 21548
rect 30331 21508 32864 21536
rect 30331 21505 30343 21508
rect 30285 21499 30343 21505
rect 32858 21496 32864 21508
rect 32916 21496 32922 21548
rect 36262 21536 36268 21548
rect 36223 21508 36268 21536
rect 36262 21496 36268 21508
rect 36320 21496 36326 21548
rect 26786 21428 26792 21480
rect 26844 21468 26850 21480
rect 28077 21471 28135 21477
rect 28077 21468 28089 21471
rect 26844 21440 28089 21468
rect 26844 21428 26850 21440
rect 28077 21437 28089 21440
rect 28123 21437 28135 21471
rect 28077 21431 28135 21437
rect 28169 21471 28227 21477
rect 28169 21437 28181 21471
rect 28215 21468 28227 21471
rect 28215 21440 29684 21468
rect 28215 21437 28227 21440
rect 28169 21431 28227 21437
rect 28092 21400 28120 21431
rect 28092 21372 29224 21400
rect 27065 21335 27123 21341
rect 27065 21301 27077 21335
rect 27111 21332 27123 21335
rect 27154 21332 27160 21344
rect 27111 21304 27160 21332
rect 27111 21301 27123 21304
rect 27065 21295 27123 21301
rect 27154 21292 27160 21304
rect 27212 21292 27218 21344
rect 29196 21341 29224 21372
rect 29656 21344 29684 21440
rect 30190 21428 30196 21480
rect 30248 21468 30254 21480
rect 31389 21471 31447 21477
rect 31389 21468 31401 21471
rect 30248 21440 31401 21468
rect 30248 21428 30254 21440
rect 31389 21437 31401 21440
rect 31435 21437 31447 21471
rect 31389 21431 31447 21437
rect 31478 21428 31484 21480
rect 31536 21468 31542 21480
rect 36081 21471 36139 21477
rect 36081 21468 36093 21471
rect 31536 21440 36093 21468
rect 31536 21428 31542 21440
rect 36081 21437 36093 21440
rect 36127 21468 36139 21471
rect 36446 21468 36452 21480
rect 36127 21440 36452 21468
rect 36127 21437 36139 21440
rect 36081 21431 36139 21437
rect 36446 21428 36452 21440
rect 36504 21428 36510 21480
rect 29181 21335 29239 21341
rect 29181 21301 29193 21335
rect 29227 21332 29239 21335
rect 29362 21332 29368 21344
rect 29227 21304 29368 21332
rect 29227 21301 29239 21304
rect 29181 21295 29239 21301
rect 29362 21292 29368 21304
rect 29420 21292 29426 21344
rect 29638 21332 29644 21344
rect 29599 21304 29644 21332
rect 29638 21292 29644 21304
rect 29696 21292 29702 21344
rect 32766 21292 32772 21344
rect 32824 21332 32830 21344
rect 34241 21335 34299 21341
rect 34241 21332 34253 21335
rect 32824 21304 34253 21332
rect 32824 21292 32830 21304
rect 34241 21301 34253 21304
rect 34287 21301 34299 21335
rect 34241 21295 34299 21301
rect 35434 21292 35440 21344
rect 35492 21332 35498 21344
rect 35529 21335 35587 21341
rect 35529 21332 35541 21335
rect 35492 21304 35541 21332
rect 35492 21292 35498 21304
rect 35529 21301 35541 21304
rect 35575 21301 35587 21335
rect 35529 21295 35587 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 27246 21128 27252 21140
rect 27207 21100 27252 21128
rect 27246 21088 27252 21100
rect 27304 21088 27310 21140
rect 27982 21128 27988 21140
rect 27943 21100 27988 21128
rect 27982 21088 27988 21100
rect 28040 21088 28046 21140
rect 29733 21131 29791 21137
rect 29733 21097 29745 21131
rect 29779 21128 29791 21131
rect 30006 21128 30012 21140
rect 29779 21100 30012 21128
rect 29779 21097 29791 21100
rect 29733 21091 29791 21097
rect 30006 21088 30012 21100
rect 30064 21088 30070 21140
rect 30926 21128 30932 21140
rect 30887 21100 30932 21128
rect 30926 21088 30932 21100
rect 30984 21088 30990 21140
rect 35526 21088 35532 21140
rect 35584 21128 35590 21140
rect 35713 21131 35771 21137
rect 35713 21128 35725 21131
rect 35584 21100 35725 21128
rect 35584 21088 35590 21100
rect 35713 21097 35725 21100
rect 35759 21097 35771 21131
rect 35713 21091 35771 21097
rect 36722 21088 36728 21140
rect 36780 21128 36786 21140
rect 36909 21131 36967 21137
rect 36909 21128 36921 21131
rect 36780 21100 36921 21128
rect 36780 21088 36786 21100
rect 36909 21097 36921 21100
rect 36955 21097 36967 21131
rect 36909 21091 36967 21097
rect 29362 21020 29368 21072
rect 29420 21060 29426 21072
rect 35894 21060 35900 21072
rect 29420 21032 35900 21060
rect 29420 21020 29426 21032
rect 35894 21020 35900 21032
rect 35952 21060 35958 21072
rect 36814 21060 36820 21072
rect 35952 21032 36820 21060
rect 35952 21020 35958 21032
rect 36814 21020 36820 21032
rect 36872 21020 36878 21072
rect 22094 20952 22100 21004
rect 22152 20992 22158 21004
rect 28537 20995 28595 21001
rect 28537 20992 28549 20995
rect 22152 20964 28549 20992
rect 22152 20952 22158 20964
rect 28537 20961 28549 20964
rect 28583 20992 28595 20995
rect 30190 20992 30196 21004
rect 28583 20964 30196 20992
rect 28583 20961 28595 20964
rect 28537 20955 28595 20961
rect 30190 20952 30196 20964
rect 30248 20992 30254 21004
rect 30285 20995 30343 21001
rect 30285 20992 30297 20995
rect 30248 20964 30297 20992
rect 30248 20952 30254 20964
rect 30285 20961 30297 20964
rect 30331 20992 30343 20995
rect 31481 20995 31539 21001
rect 31481 20992 31493 20995
rect 30331 20964 31493 20992
rect 30331 20961 30343 20964
rect 30285 20955 30343 20961
rect 31481 20961 31493 20964
rect 31527 20961 31539 20995
rect 31481 20955 31539 20961
rect 35802 20952 35808 21004
rect 35860 20992 35866 21004
rect 36265 20995 36323 21001
rect 36265 20992 36277 20995
rect 35860 20964 36277 20992
rect 35860 20952 35866 20964
rect 36265 20961 36277 20964
rect 36311 20961 36323 20995
rect 36265 20955 36323 20961
rect 29454 20884 29460 20936
rect 29512 20924 29518 20936
rect 30098 20924 30104 20936
rect 29512 20896 30104 20924
rect 29512 20884 29518 20896
rect 30098 20884 30104 20896
rect 30156 20884 30162 20936
rect 31294 20924 31300 20936
rect 31255 20896 31300 20924
rect 31294 20884 31300 20896
rect 31352 20884 31358 20936
rect 36081 20927 36139 20933
rect 36081 20893 36093 20927
rect 36127 20924 36139 20927
rect 36722 20924 36728 20936
rect 36127 20896 36728 20924
rect 36127 20893 36139 20896
rect 36081 20887 36139 20893
rect 36722 20884 36728 20896
rect 36780 20884 36786 20936
rect 28350 20856 28356 20868
rect 28263 20828 28356 20856
rect 28350 20816 28356 20828
rect 28408 20856 28414 20868
rect 31662 20856 31668 20868
rect 28408 20828 31668 20856
rect 28408 20816 28414 20828
rect 31662 20816 31668 20828
rect 31720 20816 31726 20868
rect 35253 20859 35311 20865
rect 35253 20825 35265 20859
rect 35299 20856 35311 20859
rect 35802 20856 35808 20868
rect 35299 20828 35808 20856
rect 35299 20825 35311 20828
rect 35253 20819 35311 20825
rect 35802 20816 35808 20828
rect 35860 20856 35866 20868
rect 36173 20859 36231 20865
rect 36173 20856 36185 20859
rect 35860 20828 36185 20856
rect 35860 20816 35866 20828
rect 36173 20825 36185 20828
rect 36219 20825 36231 20859
rect 36173 20819 36231 20825
rect 20990 20788 20996 20800
rect 20951 20760 20996 20788
rect 20990 20748 20996 20760
rect 21048 20748 21054 20800
rect 28445 20791 28503 20797
rect 28445 20757 28457 20791
rect 28491 20788 28503 20791
rect 28810 20788 28816 20800
rect 28491 20760 28816 20788
rect 28491 20757 28503 20760
rect 28445 20751 28503 20757
rect 28810 20748 28816 20760
rect 28868 20748 28874 20800
rect 30193 20791 30251 20797
rect 30193 20757 30205 20791
rect 30239 20788 30251 20791
rect 30742 20788 30748 20800
rect 30239 20760 30748 20788
rect 30239 20757 30251 20760
rect 30193 20751 30251 20757
rect 30742 20748 30748 20760
rect 30800 20748 30806 20800
rect 31389 20791 31447 20797
rect 31389 20757 31401 20791
rect 31435 20788 31447 20791
rect 32217 20791 32275 20797
rect 32217 20788 32229 20791
rect 31435 20760 32229 20788
rect 31435 20757 31447 20760
rect 31389 20751 31447 20757
rect 32217 20757 32229 20760
rect 32263 20788 32275 20791
rect 32306 20788 32312 20800
rect 32263 20760 32312 20788
rect 32263 20757 32275 20760
rect 32217 20751 32275 20757
rect 32306 20748 32312 20760
rect 32364 20748 32370 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 20441 20587 20499 20593
rect 20441 20553 20453 20587
rect 20487 20584 20499 20587
rect 20990 20584 20996 20596
rect 20487 20556 20996 20584
rect 20487 20553 20499 20556
rect 20441 20547 20499 20553
rect 20990 20544 20996 20556
rect 21048 20584 21054 20596
rect 27062 20584 27068 20596
rect 21048 20556 27068 20584
rect 21048 20544 21054 20556
rect 27062 20544 27068 20556
rect 27120 20544 27126 20596
rect 28350 20584 28356 20596
rect 28311 20556 28356 20584
rect 28350 20544 28356 20556
rect 28408 20544 28414 20596
rect 29549 20587 29607 20593
rect 29549 20553 29561 20587
rect 29595 20584 29607 20587
rect 29822 20584 29828 20596
rect 29595 20556 29828 20584
rect 29595 20553 29607 20556
rect 29549 20547 29607 20553
rect 29822 20544 29828 20556
rect 29880 20544 29886 20596
rect 30098 20544 30104 20596
rect 30156 20584 30162 20596
rect 31297 20587 31355 20593
rect 31297 20584 31309 20587
rect 30156 20556 31309 20584
rect 30156 20544 30162 20556
rect 31297 20553 31309 20556
rect 31343 20553 31355 20587
rect 31297 20547 31355 20553
rect 23290 20516 23296 20528
rect 22066 20488 23296 20516
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20448 20591 20451
rect 21821 20451 21879 20457
rect 21821 20448 21833 20451
rect 20579 20420 21833 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 21821 20417 21833 20420
rect 21867 20448 21879 20451
rect 22066 20448 22094 20488
rect 23290 20476 23296 20488
rect 23348 20476 23354 20528
rect 29914 20448 29920 20460
rect 21867 20420 22094 20448
rect 29875 20420 29920 20448
rect 21867 20417 21879 20420
rect 21821 20411 21879 20417
rect 29914 20408 29920 20420
rect 29972 20408 29978 20460
rect 20717 20383 20775 20389
rect 20717 20349 20729 20383
rect 20763 20380 20775 20383
rect 22094 20380 22100 20392
rect 20763 20352 22100 20380
rect 20763 20349 20775 20352
rect 20717 20343 20775 20349
rect 22094 20340 22100 20352
rect 22152 20340 22158 20392
rect 30006 20380 30012 20392
rect 29967 20352 30012 20380
rect 30006 20340 30012 20352
rect 30064 20340 30070 20392
rect 30190 20380 30196 20392
rect 30151 20352 30196 20380
rect 30190 20340 30196 20352
rect 30248 20340 30254 20392
rect 20073 20247 20131 20253
rect 20073 20213 20085 20247
rect 20119 20244 20131 20247
rect 20162 20244 20168 20256
rect 20119 20216 20168 20244
rect 20119 20213 20131 20216
rect 20073 20207 20131 20213
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 28810 20244 28816 20256
rect 28771 20216 28816 20244
rect 28810 20204 28816 20216
rect 28868 20204 28874 20256
rect 30742 20244 30748 20256
rect 30703 20216 30748 20244
rect 30742 20204 30748 20216
rect 30800 20204 30806 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 21174 20000 21180 20052
rect 21232 20040 21238 20052
rect 21358 20040 21364 20052
rect 21232 20012 21364 20040
rect 21232 20000 21238 20012
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 22833 20043 22891 20049
rect 22833 20009 22845 20043
rect 22879 20040 22891 20043
rect 22922 20040 22928 20052
rect 22879 20012 22928 20040
rect 22879 20009 22891 20012
rect 22833 20003 22891 20009
rect 20438 19904 20444 19916
rect 20399 19876 20444 19904
rect 20438 19864 20444 19876
rect 20496 19864 20502 19916
rect 21177 19907 21235 19913
rect 21177 19873 21189 19907
rect 21223 19904 21235 19907
rect 22094 19904 22100 19916
rect 21223 19876 22100 19904
rect 21223 19873 21235 19876
rect 21177 19867 21235 19873
rect 22094 19864 22100 19876
rect 22152 19864 22158 19916
rect 21269 19839 21327 19845
rect 21269 19805 21281 19839
rect 21315 19836 21327 19839
rect 22848 19836 22876 20003
rect 22922 20000 22928 20012
rect 22980 20000 22986 20052
rect 28997 20043 29055 20049
rect 28997 20009 29009 20043
rect 29043 20040 29055 20043
rect 29178 20040 29184 20052
rect 29043 20012 29184 20040
rect 29043 20009 29055 20012
rect 28997 20003 29055 20009
rect 29178 20000 29184 20012
rect 29236 20000 29242 20052
rect 29914 20000 29920 20052
rect 29972 20040 29978 20052
rect 30469 20043 30527 20049
rect 30469 20040 30481 20043
rect 29972 20012 30481 20040
rect 29972 20000 29978 20012
rect 30469 20009 30481 20012
rect 30515 20040 30527 20043
rect 32214 20040 32220 20052
rect 30515 20012 32220 20040
rect 30515 20009 30527 20012
rect 30469 20003 30527 20009
rect 32214 20000 32220 20012
rect 32272 20000 32278 20052
rect 36081 20043 36139 20049
rect 36081 20009 36093 20043
rect 36127 20040 36139 20043
rect 36262 20040 36268 20052
rect 36127 20012 36268 20040
rect 36127 20009 36139 20012
rect 36081 20003 36139 20009
rect 36262 20000 36268 20012
rect 36320 20000 36326 20052
rect 29196 19904 29224 20000
rect 29549 19907 29607 19913
rect 29549 19904 29561 19907
rect 29196 19876 29561 19904
rect 29549 19873 29561 19876
rect 29595 19873 29607 19907
rect 29549 19867 29607 19873
rect 35621 19907 35679 19913
rect 35621 19873 35633 19907
rect 35667 19904 35679 19907
rect 35894 19904 35900 19916
rect 35667 19876 35900 19904
rect 35667 19873 35679 19876
rect 35621 19867 35679 19873
rect 35894 19864 35900 19876
rect 35952 19904 35958 19916
rect 36633 19907 36691 19913
rect 36633 19904 36645 19907
rect 35952 19876 36645 19904
rect 35952 19864 35958 19876
rect 36633 19873 36645 19876
rect 36679 19873 36691 19907
rect 36633 19867 36691 19873
rect 21315 19808 22876 19836
rect 29733 19839 29791 19845
rect 21315 19805 21327 19808
rect 21269 19799 21327 19805
rect 29733 19805 29745 19839
rect 29779 19836 29791 19839
rect 29914 19836 29920 19848
rect 29779 19808 29920 19836
rect 29779 19805 29791 19808
rect 29733 19799 29791 19805
rect 29914 19796 29920 19808
rect 29972 19796 29978 19848
rect 36446 19836 36452 19848
rect 36407 19808 36452 19836
rect 36446 19796 36452 19808
rect 36504 19796 36510 19848
rect 20165 19771 20223 19777
rect 20165 19737 20177 19771
rect 20211 19768 20223 19771
rect 22281 19771 22339 19777
rect 22281 19768 22293 19771
rect 20211 19740 22293 19768
rect 20211 19737 20223 19740
rect 20165 19731 20223 19737
rect 22281 19737 22293 19740
rect 22327 19768 22339 19771
rect 30558 19768 30564 19780
rect 22327 19740 30564 19768
rect 22327 19737 22339 19740
rect 22281 19731 22339 19737
rect 30558 19728 30564 19740
rect 30616 19728 30622 19780
rect 19797 19703 19855 19709
rect 19797 19669 19809 19703
rect 19843 19700 19855 19703
rect 20070 19700 20076 19712
rect 19843 19672 20076 19700
rect 19843 19669 19855 19672
rect 19797 19663 19855 19669
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 20257 19703 20315 19709
rect 20257 19669 20269 19703
rect 20303 19700 20315 19703
rect 21174 19700 21180 19712
rect 20303 19672 21180 19700
rect 20303 19669 20315 19672
rect 20257 19663 20315 19669
rect 21174 19660 21180 19672
rect 21232 19660 21238 19712
rect 21358 19700 21364 19712
rect 21319 19672 21364 19700
rect 21358 19660 21364 19672
rect 21416 19660 21422 19712
rect 21729 19703 21787 19709
rect 21729 19669 21741 19703
rect 21775 19700 21787 19703
rect 22002 19700 22008 19712
rect 21775 19672 22008 19700
rect 21775 19669 21787 19672
rect 21729 19663 21787 19669
rect 22002 19660 22008 19672
rect 22060 19660 22066 19712
rect 29917 19703 29975 19709
rect 29917 19669 29929 19703
rect 29963 19700 29975 19703
rect 30098 19700 30104 19712
rect 29963 19672 30104 19700
rect 29963 19669 29975 19672
rect 29917 19663 29975 19669
rect 30098 19660 30104 19672
rect 30156 19660 30162 19712
rect 36541 19703 36599 19709
rect 36541 19669 36553 19703
rect 36587 19700 36599 19703
rect 37458 19700 37464 19712
rect 36587 19672 37464 19700
rect 36587 19669 36599 19672
rect 36541 19663 36599 19669
rect 37458 19660 37464 19672
rect 37516 19660 37522 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 20438 19496 20444 19508
rect 20399 19468 20444 19496
rect 20438 19456 20444 19468
rect 20496 19456 20502 19508
rect 21358 19456 21364 19508
rect 21416 19496 21422 19508
rect 21818 19496 21824 19508
rect 21416 19468 21824 19496
rect 21416 19456 21422 19468
rect 21818 19456 21824 19468
rect 21876 19456 21882 19508
rect 30285 19499 30343 19505
rect 30285 19465 30297 19499
rect 30331 19496 30343 19499
rect 32674 19496 32680 19508
rect 30331 19468 32680 19496
rect 30331 19465 30343 19468
rect 30285 19459 30343 19465
rect 32674 19456 32680 19468
rect 32732 19456 32738 19508
rect 35529 19499 35587 19505
rect 35529 19465 35541 19499
rect 35575 19465 35587 19499
rect 35529 19459 35587 19465
rect 35897 19499 35955 19505
rect 35897 19465 35909 19499
rect 35943 19496 35955 19499
rect 36078 19496 36084 19508
rect 35943 19468 36084 19496
rect 35943 19465 35955 19468
rect 35897 19459 35955 19465
rect 30650 19388 30656 19440
rect 30708 19428 30714 19440
rect 35544 19428 35572 19459
rect 36078 19456 36084 19468
rect 36136 19456 36142 19508
rect 30708 19400 35572 19428
rect 30708 19388 30714 19400
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19360 20591 19363
rect 22094 19360 22100 19372
rect 20579 19332 22100 19360
rect 20579 19329 20591 19332
rect 20533 19323 20591 19329
rect 22094 19320 22100 19332
rect 22152 19320 22158 19372
rect 30098 19360 30104 19372
rect 30059 19332 30104 19360
rect 30098 19320 30104 19332
rect 30156 19320 30162 19372
rect 35894 19360 35900 19372
rect 35820 19332 35900 19360
rect 21174 19292 21180 19304
rect 21135 19264 21180 19292
rect 21174 19252 21180 19264
rect 21232 19252 21238 19304
rect 27154 19252 27160 19304
rect 27212 19292 27218 19304
rect 33502 19292 33508 19304
rect 27212 19264 33508 19292
rect 27212 19252 27218 19264
rect 33502 19252 33508 19264
rect 33560 19252 33566 19304
rect 21818 19116 21824 19168
rect 21876 19156 21882 19168
rect 29178 19156 29184 19168
rect 21876 19128 29184 19156
rect 21876 19116 21882 19128
rect 29178 19116 29184 19128
rect 29236 19116 29242 19168
rect 29457 19159 29515 19165
rect 29457 19125 29469 19159
rect 29503 19156 29515 19159
rect 29914 19156 29920 19168
rect 29503 19128 29920 19156
rect 29503 19125 29515 19128
rect 29457 19119 29515 19125
rect 29914 19116 29920 19128
rect 29972 19116 29978 19168
rect 35069 19159 35127 19165
rect 35069 19125 35081 19159
rect 35115 19156 35127 19159
rect 35687 19159 35745 19165
rect 35687 19156 35699 19159
rect 35115 19128 35699 19156
rect 35115 19125 35127 19128
rect 35069 19119 35127 19125
rect 35687 19125 35699 19128
rect 35733 19156 35745 19159
rect 35820 19156 35848 19332
rect 35894 19320 35900 19332
rect 35952 19320 35958 19372
rect 35989 19295 36047 19301
rect 35989 19261 36001 19295
rect 36035 19292 36047 19295
rect 36538 19292 36544 19304
rect 36035 19264 36544 19292
rect 36035 19261 36047 19264
rect 35989 19255 36047 19261
rect 36538 19252 36544 19264
rect 36596 19252 36602 19304
rect 35733 19128 35848 19156
rect 35733 19125 35745 19128
rect 35687 19119 35745 19125
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 23569 18955 23627 18961
rect 23569 18921 23581 18955
rect 23615 18952 23627 18955
rect 25406 18952 25412 18964
rect 23615 18924 25412 18952
rect 23615 18921 23627 18924
rect 23569 18915 23627 18921
rect 22094 18776 22100 18828
rect 22152 18816 22158 18828
rect 22373 18819 22431 18825
rect 22373 18816 22385 18819
rect 22152 18788 22385 18816
rect 22152 18776 22158 18788
rect 22373 18785 22385 18788
rect 22419 18816 22431 18819
rect 23382 18816 23388 18828
rect 22419 18788 23388 18816
rect 22419 18785 22431 18788
rect 22373 18779 22431 18785
rect 23382 18776 23388 18788
rect 23440 18776 23446 18828
rect 22189 18751 22247 18757
rect 22189 18717 22201 18751
rect 22235 18748 22247 18751
rect 23584 18748 23612 18915
rect 25406 18912 25412 18924
rect 25464 18912 25470 18964
rect 36078 18912 36084 18964
rect 36136 18952 36142 18964
rect 36357 18955 36415 18961
rect 36357 18952 36369 18955
rect 36136 18924 36369 18952
rect 36136 18912 36142 18924
rect 36357 18921 36369 18924
rect 36403 18921 36415 18955
rect 36357 18915 36415 18921
rect 22235 18720 23612 18748
rect 22235 18717 22247 18720
rect 22189 18711 22247 18717
rect 22097 18683 22155 18689
rect 22097 18649 22109 18683
rect 22143 18680 22155 18683
rect 23017 18683 23075 18689
rect 23017 18680 23029 18683
rect 22143 18652 23029 18680
rect 22143 18649 22155 18652
rect 22097 18643 22155 18649
rect 23017 18649 23029 18652
rect 23063 18680 23075 18683
rect 26234 18680 26240 18692
rect 23063 18652 26240 18680
rect 23063 18649 23075 18652
rect 23017 18643 23075 18649
rect 26234 18640 26240 18652
rect 26292 18640 26298 18692
rect 20714 18572 20720 18624
rect 20772 18612 20778 18624
rect 21729 18615 21787 18621
rect 21729 18612 21741 18615
rect 20772 18584 21741 18612
rect 20772 18572 20778 18584
rect 21729 18581 21741 18584
rect 21775 18581 21787 18615
rect 21729 18575 21787 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 17681 18411 17739 18417
rect 17681 18377 17693 18411
rect 17727 18408 17739 18411
rect 18509 18411 18567 18417
rect 18509 18408 18521 18411
rect 17727 18380 18521 18408
rect 17727 18377 17739 18380
rect 17681 18371 17739 18377
rect 18509 18377 18521 18380
rect 18555 18408 18567 18411
rect 21082 18408 21088 18420
rect 18555 18380 21088 18408
rect 18555 18377 18567 18380
rect 18509 18371 18567 18377
rect 21082 18368 21088 18380
rect 21140 18368 21146 18420
rect 33778 18408 33784 18420
rect 33739 18380 33784 18408
rect 33778 18368 33784 18380
rect 33836 18368 33842 18420
rect 34241 18411 34299 18417
rect 34241 18377 34253 18411
rect 34287 18377 34299 18411
rect 34241 18371 34299 18377
rect 16482 18232 16488 18284
rect 16540 18272 16546 18284
rect 17589 18275 17647 18281
rect 17589 18272 17601 18275
rect 16540 18244 17601 18272
rect 16540 18232 16546 18244
rect 17589 18241 17601 18244
rect 17635 18241 17647 18275
rect 17589 18235 17647 18241
rect 33873 18275 33931 18281
rect 33873 18241 33885 18275
rect 33919 18241 33931 18275
rect 34256 18272 34284 18371
rect 34701 18275 34759 18281
rect 34701 18272 34713 18275
rect 34256 18244 34713 18272
rect 33873 18235 33931 18241
rect 34701 18241 34713 18244
rect 34747 18241 34759 18275
rect 34701 18235 34759 18241
rect 17865 18207 17923 18213
rect 17865 18173 17877 18207
rect 17911 18204 17923 18207
rect 20438 18204 20444 18216
rect 17911 18176 20444 18204
rect 17911 18173 17923 18176
rect 17865 18167 17923 18173
rect 20438 18164 20444 18176
rect 20496 18164 20502 18216
rect 33597 18207 33655 18213
rect 33597 18204 33609 18207
rect 33244 18176 33609 18204
rect 33244 18080 33272 18176
rect 33597 18173 33609 18176
rect 33643 18173 33655 18207
rect 33888 18204 33916 18235
rect 34606 18204 34612 18216
rect 33888 18176 34612 18204
rect 33597 18167 33655 18173
rect 34606 18164 34612 18176
rect 34664 18164 34670 18216
rect 15930 18028 15936 18080
rect 15988 18068 15994 18080
rect 17221 18071 17279 18077
rect 17221 18068 17233 18071
rect 15988 18040 17233 18068
rect 15988 18028 15994 18040
rect 17221 18037 17233 18040
rect 17267 18037 17279 18071
rect 17221 18031 17279 18037
rect 33045 18071 33103 18077
rect 33045 18037 33057 18071
rect 33091 18068 33103 18071
rect 33226 18068 33232 18080
rect 33091 18040 33232 18068
rect 33091 18037 33103 18040
rect 33045 18031 33103 18037
rect 33226 18028 33232 18040
rect 33284 18028 33290 18080
rect 34790 18028 34796 18080
rect 34848 18068 34854 18080
rect 34885 18071 34943 18077
rect 34885 18068 34897 18071
rect 34848 18040 34897 18068
rect 34848 18028 34854 18040
rect 34885 18037 34897 18040
rect 34931 18037 34943 18071
rect 34885 18031 34943 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 34606 17824 34612 17876
rect 34664 17864 34670 17876
rect 34701 17867 34759 17873
rect 34701 17864 34713 17867
rect 34664 17836 34713 17864
rect 34664 17824 34670 17836
rect 34701 17833 34713 17836
rect 34747 17833 34759 17867
rect 34701 17827 34759 17833
rect 16482 17484 16488 17536
rect 16540 17524 16546 17536
rect 18049 17527 18107 17533
rect 18049 17524 18061 17527
rect 16540 17496 18061 17524
rect 16540 17484 16546 17496
rect 18049 17493 18061 17496
rect 18095 17493 18107 17527
rect 18049 17487 18107 17493
rect 34606 17484 34612 17536
rect 34664 17524 34670 17536
rect 37734 17524 37740 17536
rect 34664 17496 37740 17524
rect 34664 17484 34670 17496
rect 37734 17484 37740 17496
rect 37792 17484 37798 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 16942 17280 16948 17332
rect 17000 17320 17006 17332
rect 17494 17320 17500 17332
rect 17000 17292 17500 17320
rect 17000 17280 17006 17292
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 18414 17280 18420 17332
rect 18472 17320 18478 17332
rect 19061 17323 19119 17329
rect 19061 17320 19073 17323
rect 18472 17292 19073 17320
rect 18472 17280 18478 17292
rect 19061 17289 19073 17292
rect 19107 17320 19119 17323
rect 21542 17320 21548 17332
rect 19107 17292 21548 17320
rect 19107 17289 19119 17292
rect 19061 17283 19119 17289
rect 21542 17280 21548 17292
rect 21600 17280 21606 17332
rect 27065 17323 27123 17329
rect 27065 17320 27077 17323
rect 26206 17292 27077 17320
rect 25501 17187 25559 17193
rect 25501 17184 25513 17187
rect 25332 17156 25513 17184
rect 25130 17076 25136 17128
rect 25188 17116 25194 17128
rect 25225 17119 25283 17125
rect 25225 17116 25237 17119
rect 25188 17088 25237 17116
rect 25188 17076 25194 17088
rect 25225 17085 25237 17088
rect 25271 17085 25283 17119
rect 25225 17079 25283 17085
rect 18322 17008 18328 17060
rect 18380 17048 18386 17060
rect 19521 17051 19579 17057
rect 19521 17048 19533 17051
rect 18380 17020 19533 17048
rect 18380 17008 18386 17020
rect 19521 17017 19533 17020
rect 19567 17017 19579 17051
rect 19521 17011 19579 17017
rect 25332 16980 25360 17156
rect 25501 17153 25513 17156
rect 25547 17153 25559 17187
rect 25501 17147 25559 17153
rect 25409 17119 25467 17125
rect 25409 17085 25421 17119
rect 25455 17116 25467 17119
rect 26206 17116 26234 17292
rect 27065 17289 27077 17292
rect 27111 17320 27123 17323
rect 33962 17320 33968 17332
rect 27111 17292 33968 17320
rect 27111 17289 27123 17292
rect 27065 17283 27123 17289
rect 33962 17280 33968 17292
rect 34020 17280 34026 17332
rect 25455 17088 26234 17116
rect 25455 17085 25467 17088
rect 25409 17079 25467 17085
rect 25869 17051 25927 17057
rect 25869 17017 25881 17051
rect 25915 17048 25927 17051
rect 26418 17048 26424 17060
rect 25915 17020 26424 17048
rect 25915 17017 25927 17020
rect 25869 17011 25927 17017
rect 26418 17008 26424 17020
rect 26476 17008 26482 17060
rect 29730 17048 29736 17060
rect 26896 17020 29736 17048
rect 26329 16983 26387 16989
rect 26329 16980 26341 16983
rect 25332 16952 26341 16980
rect 26329 16949 26341 16952
rect 26375 16980 26387 16983
rect 26896 16980 26924 17020
rect 29730 17008 29736 17020
rect 29788 17008 29794 17060
rect 26375 16952 26924 16980
rect 26375 16949 26387 16952
rect 26329 16943 26387 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 22373 16779 22431 16785
rect 22373 16745 22385 16779
rect 22419 16776 22431 16779
rect 24394 16776 24400 16788
rect 22419 16748 24400 16776
rect 22419 16745 22431 16748
rect 22373 16739 22431 16745
rect 22388 16708 22416 16739
rect 24394 16736 24400 16748
rect 24452 16736 24458 16788
rect 21008 16680 22416 16708
rect 18414 16640 18420 16652
rect 18375 16612 18420 16640
rect 18414 16600 18420 16612
rect 18472 16600 18478 16652
rect 18601 16643 18659 16649
rect 18601 16609 18613 16643
rect 18647 16640 18659 16643
rect 18966 16640 18972 16652
rect 18647 16612 18972 16640
rect 18647 16609 18659 16612
rect 18601 16603 18659 16609
rect 18966 16600 18972 16612
rect 19024 16640 19030 16652
rect 20438 16640 20444 16652
rect 19024 16612 20444 16640
rect 19024 16600 19030 16612
rect 20438 16600 20444 16612
rect 20496 16640 20502 16652
rect 21008 16649 21036 16680
rect 20993 16643 21051 16649
rect 20496 16612 20944 16640
rect 20496 16600 20502 16612
rect 20916 16572 20944 16612
rect 20993 16609 21005 16643
rect 21039 16609 21051 16643
rect 20993 16603 21051 16609
rect 21085 16643 21143 16649
rect 21085 16609 21097 16643
rect 21131 16609 21143 16643
rect 21085 16603 21143 16609
rect 21100 16572 21128 16603
rect 20916 16544 21128 16572
rect 23382 16532 23388 16584
rect 23440 16572 23446 16584
rect 25130 16572 25136 16584
rect 23440 16544 25136 16572
rect 23440 16532 23446 16544
rect 25130 16532 25136 16544
rect 25188 16532 25194 16584
rect 19334 16464 19340 16516
rect 19392 16504 19398 16516
rect 19705 16507 19763 16513
rect 19705 16504 19717 16507
rect 19392 16476 19717 16504
rect 19392 16464 19398 16476
rect 19705 16473 19717 16476
rect 19751 16504 19763 16507
rect 22738 16504 22744 16516
rect 19751 16476 22744 16504
rect 19751 16473 19763 16476
rect 19705 16467 19763 16473
rect 22738 16464 22744 16476
rect 22796 16464 22802 16516
rect 16850 16396 16856 16448
rect 16908 16436 16914 16448
rect 17957 16439 18015 16445
rect 17957 16436 17969 16439
rect 16908 16408 17969 16436
rect 16908 16396 16914 16408
rect 17957 16405 17969 16408
rect 18003 16405 18015 16439
rect 18322 16436 18328 16448
rect 18283 16408 18328 16436
rect 17957 16399 18015 16405
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 18506 16396 18512 16448
rect 18564 16436 18570 16448
rect 20533 16439 20591 16445
rect 20533 16436 20545 16439
rect 18564 16408 20545 16436
rect 18564 16396 18570 16408
rect 20533 16405 20545 16408
rect 20579 16405 20591 16439
rect 20533 16399 20591 16405
rect 20901 16439 20959 16445
rect 20901 16405 20913 16439
rect 20947 16436 20959 16439
rect 21729 16439 21787 16445
rect 21729 16436 21741 16439
rect 20947 16408 21741 16436
rect 20947 16405 20959 16408
rect 20901 16399 20959 16405
rect 21729 16405 21741 16408
rect 21775 16436 21787 16439
rect 21818 16436 21824 16448
rect 21775 16408 21824 16436
rect 21775 16405 21787 16408
rect 21729 16399 21787 16405
rect 21818 16396 21824 16408
rect 21876 16396 21882 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 17405 16235 17463 16241
rect 17405 16201 17417 16235
rect 17451 16232 17463 16235
rect 17954 16232 17960 16244
rect 17451 16204 17960 16232
rect 17451 16201 17463 16204
rect 17405 16195 17463 16201
rect 17954 16192 17960 16204
rect 18012 16232 18018 16244
rect 18598 16232 18604 16244
rect 18012 16204 18604 16232
rect 18012 16192 18018 16204
rect 18598 16192 18604 16204
rect 18656 16192 18662 16244
rect 19153 16235 19211 16241
rect 19153 16201 19165 16235
rect 19199 16232 19211 16235
rect 19334 16232 19340 16244
rect 19199 16204 19340 16232
rect 19199 16201 19211 16204
rect 19153 16195 19211 16201
rect 19334 16192 19340 16204
rect 19392 16192 19398 16244
rect 19061 16167 19119 16173
rect 19061 16133 19073 16167
rect 19107 16164 19119 16167
rect 19426 16164 19432 16176
rect 19107 16136 19432 16164
rect 19107 16133 19119 16136
rect 19061 16127 19119 16133
rect 19426 16124 19432 16136
rect 19484 16164 19490 16176
rect 19981 16167 20039 16173
rect 19981 16164 19993 16167
rect 19484 16136 19993 16164
rect 19484 16124 19490 16136
rect 19981 16133 19993 16136
rect 20027 16133 20039 16167
rect 19981 16127 20039 16133
rect 23201 16167 23259 16173
rect 23201 16133 23213 16167
rect 23247 16164 23259 16167
rect 24026 16164 24032 16176
rect 23247 16136 24032 16164
rect 23247 16133 23259 16136
rect 23201 16127 23259 16133
rect 24026 16124 24032 16136
rect 24084 16164 24090 16176
rect 24489 16167 24547 16173
rect 24489 16164 24501 16167
rect 24084 16136 24501 16164
rect 24084 16124 24090 16136
rect 24489 16133 24501 16136
rect 24535 16133 24547 16167
rect 24489 16127 24547 16133
rect 22002 16096 22008 16108
rect 21963 16068 22008 16096
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 23109 16099 23167 16105
rect 23109 16065 23121 16099
rect 23155 16096 23167 16099
rect 23937 16099 23995 16105
rect 23937 16096 23949 16099
rect 23155 16068 23949 16096
rect 23155 16065 23167 16068
rect 23109 16059 23167 16065
rect 23937 16065 23949 16068
rect 23983 16096 23995 16099
rect 24854 16096 24860 16108
rect 23983 16068 24860 16096
rect 23983 16065 23995 16068
rect 23937 16059 23995 16065
rect 24854 16056 24860 16068
rect 24912 16056 24918 16108
rect 18966 16028 18972 16040
rect 18927 16000 18972 16028
rect 18966 15988 18972 16000
rect 19024 15988 19030 16040
rect 22189 16031 22247 16037
rect 22189 15997 22201 16031
rect 22235 16028 22247 16031
rect 22646 16028 22652 16040
rect 22235 16000 22652 16028
rect 22235 15997 22247 16000
rect 22189 15991 22247 15997
rect 22646 15988 22652 16000
rect 22704 15988 22710 16040
rect 23290 16028 23296 16040
rect 23251 16000 23296 16028
rect 23290 15988 23296 16000
rect 23348 15988 23354 16040
rect 19426 15852 19432 15904
rect 19484 15892 19490 15904
rect 19521 15895 19579 15901
rect 19521 15892 19533 15895
rect 19484 15864 19533 15892
rect 19484 15852 19490 15864
rect 19521 15861 19533 15864
rect 19567 15861 19579 15895
rect 19521 15855 19579 15861
rect 21726 15852 21732 15904
rect 21784 15892 21790 15904
rect 21821 15895 21879 15901
rect 21821 15892 21833 15895
rect 21784 15864 21833 15892
rect 21784 15852 21790 15864
rect 21821 15861 21833 15864
rect 21867 15861 21879 15895
rect 21821 15855 21879 15861
rect 22554 15852 22560 15904
rect 22612 15892 22618 15904
rect 22741 15895 22799 15901
rect 22741 15892 22753 15895
rect 22612 15864 22753 15892
rect 22612 15852 22618 15864
rect 22741 15861 22753 15864
rect 22787 15861 22799 15895
rect 22741 15855 22799 15861
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 21269 15691 21327 15697
rect 21269 15688 21281 15691
rect 20456 15660 21281 15688
rect 17954 15620 17960 15632
rect 16960 15592 17960 15620
rect 16960 15561 16988 15592
rect 17954 15580 17960 15592
rect 18012 15580 18018 15632
rect 16945 15555 17003 15561
rect 16945 15521 16957 15555
rect 16991 15521 17003 15555
rect 16945 15515 17003 15521
rect 17129 15555 17187 15561
rect 17129 15521 17141 15555
rect 17175 15552 17187 15555
rect 18966 15552 18972 15564
rect 17175 15524 18972 15552
rect 17175 15521 17187 15524
rect 17129 15515 17187 15521
rect 18966 15512 18972 15524
rect 19024 15512 19030 15564
rect 20456 15561 20484 15660
rect 21269 15657 21281 15660
rect 21315 15688 21327 15691
rect 22186 15688 22192 15700
rect 21315 15660 22192 15688
rect 21315 15657 21327 15660
rect 21269 15651 21327 15657
rect 22186 15648 22192 15660
rect 22244 15648 22250 15700
rect 24581 15691 24639 15697
rect 24581 15657 24593 15691
rect 24627 15688 24639 15691
rect 30650 15688 30656 15700
rect 24627 15660 30656 15688
rect 24627 15657 24639 15660
rect 24581 15651 24639 15657
rect 30650 15648 30656 15660
rect 30708 15648 30714 15700
rect 21913 15623 21971 15629
rect 21913 15589 21925 15623
rect 21959 15620 21971 15623
rect 25590 15620 25596 15632
rect 21959 15592 25596 15620
rect 21959 15589 21971 15592
rect 21913 15583 21971 15589
rect 25590 15580 25596 15592
rect 25648 15580 25654 15632
rect 26418 15580 26424 15632
rect 26476 15620 26482 15632
rect 26605 15623 26663 15629
rect 26476 15592 26556 15620
rect 26476 15580 26482 15592
rect 20441 15555 20499 15561
rect 20441 15521 20453 15555
rect 20487 15521 20499 15555
rect 20441 15515 20499 15521
rect 20625 15555 20683 15561
rect 20625 15521 20637 15555
rect 20671 15552 20683 15555
rect 23290 15552 23296 15564
rect 20671 15524 23296 15552
rect 20671 15521 20683 15524
rect 20625 15515 20683 15521
rect 23290 15512 23296 15524
rect 23348 15512 23354 15564
rect 17402 15444 17408 15496
rect 17460 15484 17466 15496
rect 17865 15487 17923 15493
rect 17865 15484 17877 15487
rect 17460 15456 17877 15484
rect 17460 15444 17466 15456
rect 17865 15453 17877 15456
rect 17911 15453 17923 15487
rect 17865 15447 17923 15453
rect 18049 15487 18107 15493
rect 18049 15453 18061 15487
rect 18095 15484 18107 15487
rect 20346 15484 20352 15496
rect 18095 15456 20352 15484
rect 18095 15453 18107 15456
rect 18049 15447 18107 15453
rect 20346 15444 20352 15456
rect 20404 15444 20410 15496
rect 21726 15484 21732 15496
rect 21687 15456 21732 15484
rect 21726 15444 21732 15456
rect 21784 15444 21790 15496
rect 22373 15487 22431 15493
rect 22373 15453 22385 15487
rect 22419 15453 22431 15487
rect 22554 15484 22560 15496
rect 22515 15456 22560 15484
rect 22373 15447 22431 15453
rect 16853 15419 16911 15425
rect 16853 15385 16865 15419
rect 16899 15416 16911 15419
rect 17494 15416 17500 15428
rect 16899 15388 17500 15416
rect 16899 15385 16911 15388
rect 16853 15379 16911 15385
rect 17494 15376 17500 15388
rect 17552 15376 17558 15428
rect 22388 15416 22416 15447
rect 22554 15444 22560 15456
rect 22612 15444 22618 15496
rect 22741 15487 22799 15493
rect 22741 15453 22753 15487
rect 22787 15484 22799 15487
rect 23201 15487 23259 15493
rect 23201 15484 23213 15487
rect 22787 15456 23213 15484
rect 22787 15453 22799 15456
rect 22741 15447 22799 15453
rect 23201 15453 23213 15456
rect 23247 15453 23259 15487
rect 24394 15484 24400 15496
rect 24355 15456 24400 15484
rect 23201 15447 23259 15453
rect 24394 15444 24400 15456
rect 24452 15444 24458 15496
rect 26050 15444 26056 15496
rect 26108 15484 26114 15496
rect 26237 15487 26295 15493
rect 26237 15484 26249 15487
rect 26108 15456 26249 15484
rect 26108 15444 26114 15456
rect 26237 15453 26249 15456
rect 26283 15453 26295 15487
rect 26237 15447 26295 15453
rect 26441 15487 26499 15493
rect 26441 15453 26453 15487
rect 26487 15484 26499 15487
rect 26528 15484 26556 15592
rect 26605 15589 26617 15623
rect 26651 15620 26663 15623
rect 30282 15620 30288 15632
rect 26651 15592 30288 15620
rect 26651 15589 26663 15592
rect 26605 15583 26663 15589
rect 30282 15580 30288 15592
rect 30340 15580 30346 15632
rect 36081 15555 36139 15561
rect 36081 15521 36093 15555
rect 36127 15552 36139 15555
rect 36262 15552 36268 15564
rect 36127 15524 36268 15552
rect 36127 15521 36139 15524
rect 36081 15515 36139 15521
rect 36262 15512 36268 15524
rect 36320 15552 36326 15564
rect 37093 15555 37151 15561
rect 37093 15552 37105 15555
rect 36320 15524 37105 15552
rect 36320 15512 36326 15524
rect 37093 15521 37105 15524
rect 37139 15521 37151 15555
rect 37093 15515 37151 15521
rect 26487 15456 26556 15484
rect 26487 15453 26499 15456
rect 26441 15447 26499 15453
rect 26602 15444 26608 15496
rect 26660 15484 26666 15496
rect 27801 15487 27859 15493
rect 26660 15456 27476 15484
rect 26660 15444 26666 15456
rect 22646 15416 22652 15428
rect 22388 15388 22652 15416
rect 22646 15376 22652 15388
rect 22704 15376 22710 15428
rect 23400 15388 26648 15416
rect 27448 15402 27476 15456
rect 27801 15453 27813 15487
rect 27847 15484 27859 15487
rect 28353 15487 28411 15493
rect 27847 15456 28120 15484
rect 27847 15453 27859 15456
rect 27801 15447 27859 15453
rect 28092 15416 28120 15456
rect 28353 15453 28365 15487
rect 28399 15484 28411 15487
rect 32122 15484 32128 15496
rect 28399 15456 32128 15484
rect 28399 15453 28411 15456
rect 28353 15447 28411 15453
rect 32122 15444 32128 15456
rect 32180 15444 32186 15496
rect 33134 15444 33140 15496
rect 33192 15484 33198 15496
rect 37737 15487 37795 15493
rect 37737 15484 37749 15487
rect 33192 15456 37749 15484
rect 33192 15444 33198 15456
rect 37737 15453 37749 15456
rect 37783 15453 37795 15487
rect 37737 15447 37795 15453
rect 33318 15416 33324 15428
rect 28092 15388 33324 15416
rect 15470 15308 15476 15360
rect 15528 15348 15534 15360
rect 16485 15351 16543 15357
rect 16485 15348 16497 15351
rect 15528 15320 16497 15348
rect 15528 15308 15534 15320
rect 16485 15317 16497 15320
rect 16531 15317 16543 15351
rect 16485 15311 16543 15317
rect 18233 15351 18291 15357
rect 18233 15317 18245 15351
rect 18279 15348 18291 15351
rect 19242 15348 19248 15360
rect 18279 15320 19248 15348
rect 18279 15317 18291 15320
rect 18233 15311 18291 15317
rect 19242 15308 19248 15320
rect 19300 15308 19306 15360
rect 19978 15348 19984 15360
rect 19939 15320 19984 15348
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 20349 15351 20407 15357
rect 20349 15317 20361 15351
rect 20395 15348 20407 15351
rect 20898 15348 20904 15360
rect 20395 15320 20904 15348
rect 20395 15317 20407 15320
rect 20349 15311 20407 15317
rect 20898 15308 20904 15320
rect 20956 15308 20962 15360
rect 23400 15357 23428 15388
rect 23385 15351 23443 15357
rect 23385 15317 23397 15351
rect 23431 15317 23443 15351
rect 25406 15348 25412 15360
rect 25367 15320 25412 15348
rect 23385 15311 23443 15317
rect 25406 15308 25412 15320
rect 25464 15308 25470 15360
rect 25498 15308 25504 15360
rect 25556 15348 25562 15360
rect 26510 15348 26516 15360
rect 25556 15320 26516 15348
rect 25556 15308 25562 15320
rect 26510 15308 26516 15320
rect 26568 15308 26574 15360
rect 26620 15348 26648 15388
rect 33318 15376 33324 15388
rect 33376 15376 33382 15428
rect 27522 15348 27528 15360
rect 26620 15320 27528 15348
rect 27522 15308 27528 15320
rect 27580 15308 27586 15360
rect 36446 15308 36452 15360
rect 36504 15348 36510 15360
rect 36541 15351 36599 15357
rect 36541 15348 36553 15351
rect 36504 15320 36553 15348
rect 36504 15308 36510 15320
rect 36541 15317 36553 15320
rect 36587 15317 36599 15351
rect 36906 15348 36912 15360
rect 36867 15320 36912 15348
rect 36541 15311 36599 15317
rect 36906 15308 36912 15320
rect 36964 15308 36970 15360
rect 37001 15351 37059 15357
rect 37001 15317 37013 15351
rect 37047 15348 37059 15351
rect 37366 15348 37372 15360
rect 37047 15320 37372 15348
rect 37047 15317 37059 15320
rect 37001 15311 37059 15317
rect 37366 15308 37372 15320
rect 37424 15308 37430 15360
rect 37918 15348 37924 15360
rect 37879 15320 37924 15348
rect 37918 15308 37924 15320
rect 37976 15308 37982 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 17310 15104 17316 15156
rect 17368 15144 17374 15156
rect 18325 15147 18383 15153
rect 18325 15144 18337 15147
rect 17368 15116 18337 15144
rect 17368 15104 17374 15116
rect 18325 15113 18337 15116
rect 18371 15144 18383 15147
rect 20254 15144 20260 15156
rect 18371 15116 20260 15144
rect 18371 15113 18383 15116
rect 18325 15107 18383 15113
rect 20254 15104 20260 15116
rect 20312 15104 20318 15156
rect 20346 15104 20352 15156
rect 20404 15144 20410 15156
rect 21821 15147 21879 15153
rect 21821 15144 21833 15147
rect 20404 15116 21833 15144
rect 20404 15104 20410 15116
rect 21821 15113 21833 15116
rect 21867 15113 21879 15147
rect 21821 15107 21879 15113
rect 23845 15147 23903 15153
rect 23845 15113 23857 15147
rect 23891 15144 23903 15147
rect 24394 15144 24400 15156
rect 23891 15116 24400 15144
rect 23891 15113 23903 15116
rect 23845 15107 23903 15113
rect 24394 15104 24400 15116
rect 24452 15104 24458 15156
rect 24946 15144 24952 15156
rect 24907 15116 24952 15144
rect 24946 15104 24952 15116
rect 25004 15104 25010 15156
rect 32493 15147 32551 15153
rect 32493 15113 32505 15147
rect 32539 15144 32551 15147
rect 33134 15144 33140 15156
rect 32539 15116 33140 15144
rect 32539 15113 32551 15116
rect 32493 15107 32551 15113
rect 33134 15104 33140 15116
rect 33192 15104 33198 15156
rect 19889 15079 19947 15085
rect 19889 15045 19901 15079
rect 19935 15076 19947 15079
rect 20622 15076 20628 15088
rect 19935 15048 20628 15076
rect 19935 15045 19947 15048
rect 19889 15039 19947 15045
rect 20622 15036 20628 15048
rect 20680 15036 20686 15088
rect 21634 15036 21640 15088
rect 21692 15076 21698 15088
rect 22281 15079 22339 15085
rect 22281 15076 22293 15079
rect 21692 15048 22293 15076
rect 21692 15036 21698 15048
rect 22281 15045 22293 15048
rect 22327 15045 22339 15079
rect 22281 15039 22339 15045
rect 24857 15079 24915 15085
rect 24857 15045 24869 15079
rect 24903 15076 24915 15079
rect 25406 15076 25412 15088
rect 24903 15048 25412 15076
rect 24903 15045 24915 15048
rect 24857 15039 24915 15045
rect 25406 15036 25412 15048
rect 25464 15036 25470 15088
rect 19797 15011 19855 15017
rect 19797 14977 19809 15011
rect 19843 15008 19855 15011
rect 20990 15008 20996 15020
rect 19843 14980 20996 15008
rect 19843 14977 19855 14980
rect 19797 14971 19855 14977
rect 20990 14968 20996 14980
rect 21048 14968 21054 15020
rect 22186 15008 22192 15020
rect 22147 14980 22192 15008
rect 22186 14968 22192 14980
rect 22244 14968 22250 15020
rect 23661 15011 23719 15017
rect 23661 14977 23673 15011
rect 23707 15008 23719 15011
rect 23707 14980 24532 15008
rect 23707 14977 23719 14980
rect 23661 14971 23719 14977
rect 18966 14900 18972 14952
rect 19024 14940 19030 14952
rect 19981 14943 20039 14949
rect 19981 14940 19993 14943
rect 19024 14912 19993 14940
rect 19024 14900 19030 14912
rect 19981 14909 19993 14912
rect 20027 14940 20039 14943
rect 22373 14943 22431 14949
rect 22373 14940 22385 14943
rect 20027 14912 22385 14940
rect 20027 14909 20039 14912
rect 19981 14903 20039 14909
rect 22373 14909 22385 14912
rect 22419 14909 22431 14943
rect 22373 14903 22431 14909
rect 22646 14900 22652 14952
rect 22704 14940 22710 14952
rect 23477 14943 23535 14949
rect 23477 14940 23489 14943
rect 22704 14912 23489 14940
rect 22704 14900 22710 14912
rect 23477 14909 23489 14912
rect 23523 14940 23535 14943
rect 23523 14912 23704 14940
rect 23523 14909 23535 14912
rect 23477 14903 23535 14909
rect 20898 14872 20904 14884
rect 20811 14844 20904 14872
rect 20898 14832 20904 14844
rect 20956 14872 20962 14884
rect 20956 14844 22094 14872
rect 20956 14832 20962 14844
rect 17218 14804 17224 14816
rect 17179 14776 17224 14804
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 17402 14764 17408 14816
rect 17460 14804 17466 14816
rect 17681 14807 17739 14813
rect 17681 14804 17693 14807
rect 17460 14776 17693 14804
rect 17460 14764 17466 14776
rect 17681 14773 17693 14776
rect 17727 14773 17739 14807
rect 17681 14767 17739 14773
rect 18966 14764 18972 14816
rect 19024 14804 19030 14816
rect 19429 14807 19487 14813
rect 19429 14804 19441 14807
rect 19024 14776 19441 14804
rect 19024 14764 19030 14776
rect 19429 14773 19441 14776
rect 19475 14773 19487 14807
rect 22066 14804 22094 14844
rect 23566 14804 23572 14816
rect 22066 14776 23572 14804
rect 19429 14767 19487 14773
rect 23566 14764 23572 14776
rect 23624 14764 23630 14816
rect 23676 14804 23704 14912
rect 24504 14881 24532 14980
rect 25314 14968 25320 15020
rect 25372 15008 25378 15020
rect 26237 15011 26295 15017
rect 26237 15008 26249 15011
rect 25372 14980 26249 15008
rect 25372 14968 25378 14980
rect 26237 14977 26249 14980
rect 26283 14977 26295 15011
rect 30282 15008 30288 15020
rect 30243 14980 30288 15008
rect 26237 14971 26295 14977
rect 30282 14968 30288 14980
rect 30340 14968 30346 15020
rect 32122 15008 32128 15020
rect 32083 14980 32128 15008
rect 32122 14968 32128 14980
rect 32180 14968 32186 15020
rect 32309 15011 32367 15017
rect 32309 14977 32321 15011
rect 32355 14977 32367 15011
rect 32309 14971 32367 14977
rect 25130 14940 25136 14952
rect 25091 14912 25136 14940
rect 25130 14900 25136 14912
rect 25188 14940 25194 14952
rect 25498 14940 25504 14952
rect 25188 14912 25504 14940
rect 25188 14900 25194 14912
rect 25498 14900 25504 14912
rect 25556 14900 25562 14952
rect 26050 14940 26056 14952
rect 26011 14912 26056 14940
rect 26050 14900 26056 14912
rect 26108 14900 26114 14952
rect 32324 14940 32352 14971
rect 31496 14912 32352 14940
rect 24489 14875 24547 14881
rect 24489 14841 24501 14875
rect 24535 14841 24547 14875
rect 24489 14835 24547 14841
rect 26068 14804 26096 14900
rect 29914 14832 29920 14884
rect 29972 14872 29978 14884
rect 30190 14872 30196 14884
rect 29972 14844 30196 14872
rect 29972 14832 29978 14844
rect 30190 14832 30196 14844
rect 30248 14872 30254 14884
rect 31496 14881 31524 14912
rect 31481 14875 31539 14881
rect 31481 14872 31493 14875
rect 30248 14844 31493 14872
rect 30248 14832 30254 14844
rect 31481 14841 31493 14844
rect 31527 14841 31539 14875
rect 31481 14835 31539 14841
rect 23676 14776 26096 14804
rect 26421 14807 26479 14813
rect 26421 14773 26433 14807
rect 26467 14804 26479 14807
rect 28534 14804 28540 14816
rect 26467 14776 28540 14804
rect 26467 14773 26479 14776
rect 26421 14767 26479 14773
rect 28534 14764 28540 14776
rect 28592 14764 28598 14816
rect 30466 14804 30472 14816
rect 30427 14776 30472 14804
rect 30466 14764 30472 14776
rect 30524 14764 30530 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 19150 14560 19156 14612
rect 19208 14600 19214 14612
rect 19245 14603 19303 14609
rect 19245 14600 19257 14603
rect 19208 14572 19257 14600
rect 19208 14560 19214 14572
rect 19245 14569 19257 14572
rect 19291 14569 19303 14603
rect 19245 14563 19303 14569
rect 20533 14603 20591 14609
rect 20533 14569 20545 14603
rect 20579 14600 20591 14603
rect 20622 14600 20628 14612
rect 20579 14572 20628 14600
rect 20579 14569 20591 14572
rect 20533 14563 20591 14569
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 20990 14600 20996 14612
rect 20951 14572 20996 14600
rect 20990 14560 20996 14572
rect 21048 14560 21054 14612
rect 21634 14560 21640 14612
rect 21692 14600 21698 14612
rect 22649 14603 22707 14609
rect 22649 14600 22661 14603
rect 21692 14572 22661 14600
rect 21692 14560 21698 14572
rect 22649 14569 22661 14572
rect 22695 14569 22707 14603
rect 25314 14600 25320 14612
rect 25275 14572 25320 14600
rect 22649 14563 22707 14569
rect 25314 14560 25320 14572
rect 25372 14560 25378 14612
rect 26418 14600 26424 14612
rect 26379 14572 26424 14600
rect 26418 14560 26424 14572
rect 26476 14560 26482 14612
rect 24946 14492 24952 14544
rect 25004 14532 25010 14544
rect 25777 14535 25835 14541
rect 25777 14532 25789 14535
rect 25004 14504 25789 14532
rect 25004 14492 25010 14504
rect 25777 14501 25789 14504
rect 25823 14501 25835 14535
rect 25777 14495 25835 14501
rect 17221 14467 17279 14473
rect 17221 14433 17233 14467
rect 17267 14464 17279 14467
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 17267 14436 18429 14464
rect 17267 14433 17279 14436
rect 17221 14427 17279 14433
rect 18417 14433 18429 14436
rect 18463 14464 18475 14467
rect 18874 14464 18880 14476
rect 18463 14436 18880 14464
rect 18463 14433 18475 14436
rect 18417 14427 18475 14433
rect 18874 14424 18880 14436
rect 18932 14424 18938 14476
rect 24765 14467 24823 14473
rect 24765 14433 24777 14467
rect 24811 14464 24823 14467
rect 25130 14464 25136 14476
rect 24811 14436 25136 14464
rect 24811 14433 24823 14436
rect 24765 14427 24823 14433
rect 25130 14424 25136 14436
rect 25188 14424 25194 14476
rect 25406 14424 25412 14476
rect 25464 14464 25470 14476
rect 33686 14464 33692 14476
rect 25464 14436 33692 14464
rect 25464 14424 25470 14436
rect 33686 14424 33692 14436
rect 33744 14424 33750 14476
rect 36262 14464 36268 14476
rect 35866 14436 36268 14464
rect 15289 14399 15347 14405
rect 15289 14365 15301 14399
rect 15335 14365 15347 14399
rect 15470 14396 15476 14408
rect 15431 14368 15476 14396
rect 15289 14359 15347 14365
rect 15304 14328 15332 14359
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 17034 14356 17040 14408
rect 17092 14396 17098 14408
rect 26602 14396 26608 14408
rect 17092 14368 26608 14396
rect 17092 14356 17098 14368
rect 26602 14356 26608 14368
rect 26660 14356 26666 14408
rect 28534 14396 28540 14408
rect 28495 14368 28540 14396
rect 28534 14356 28540 14368
rect 28592 14356 28598 14408
rect 32401 14399 32459 14405
rect 32401 14396 32413 14399
rect 31864 14368 32413 14396
rect 15838 14328 15844 14340
rect 15304 14300 15844 14328
rect 15838 14288 15844 14300
rect 15896 14288 15902 14340
rect 16945 14331 17003 14337
rect 16945 14297 16957 14331
rect 16991 14328 17003 14331
rect 17218 14328 17224 14340
rect 16991 14300 17224 14328
rect 16991 14297 17003 14300
rect 16945 14291 17003 14297
rect 17218 14288 17224 14300
rect 17276 14328 17282 14340
rect 19334 14328 19340 14340
rect 17276 14300 19340 14328
rect 17276 14288 17282 14300
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 24857 14331 24915 14337
rect 24857 14297 24869 14331
rect 24903 14328 24915 14331
rect 26418 14328 26424 14340
rect 24903 14300 26424 14328
rect 24903 14297 24915 14300
rect 24857 14291 24915 14297
rect 26418 14288 26424 14300
rect 26476 14288 26482 14340
rect 31864 14272 31892 14368
rect 32401 14365 32413 14368
rect 32447 14365 32459 14399
rect 32582 14396 32588 14408
rect 32543 14368 32588 14396
rect 32401 14359 32459 14365
rect 32582 14356 32588 14368
rect 32640 14356 32646 14408
rect 32769 14399 32827 14405
rect 32769 14365 32781 14399
rect 32815 14396 32827 14399
rect 33229 14399 33287 14405
rect 33229 14396 33241 14399
rect 32815 14368 33241 14396
rect 32815 14365 32827 14368
rect 32769 14359 32827 14365
rect 33229 14365 33241 14368
rect 33275 14365 33287 14399
rect 33229 14359 33287 14365
rect 15654 14260 15660 14272
rect 15615 14232 15660 14260
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 16574 14260 16580 14272
rect 16535 14232 16580 14260
rect 16574 14220 16580 14232
rect 16632 14220 16638 14272
rect 17037 14263 17095 14269
rect 17037 14229 17049 14263
rect 17083 14260 17095 14263
rect 17310 14260 17316 14272
rect 17083 14232 17316 14260
rect 17083 14229 17095 14232
rect 17037 14223 17095 14229
rect 17310 14220 17316 14232
rect 17368 14220 17374 14272
rect 17770 14260 17776 14272
rect 17731 14232 17776 14260
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 18138 14260 18144 14272
rect 18099 14232 18144 14260
rect 18138 14220 18144 14232
rect 18196 14220 18202 14272
rect 18233 14263 18291 14269
rect 18233 14229 18245 14263
rect 18279 14260 18291 14263
rect 19150 14260 19156 14272
rect 18279 14232 19156 14260
rect 18279 14229 18291 14232
rect 18233 14223 18291 14229
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 24949 14263 25007 14269
rect 24949 14229 24961 14263
rect 24995 14260 25007 14263
rect 25406 14260 25412 14272
rect 24995 14232 25412 14260
rect 24995 14229 25007 14232
rect 24949 14223 25007 14229
rect 25406 14220 25412 14232
rect 25464 14220 25470 14272
rect 28721 14263 28779 14269
rect 28721 14229 28733 14263
rect 28767 14260 28779 14263
rect 30282 14260 30288 14272
rect 28767 14232 30288 14260
rect 28767 14229 28779 14232
rect 28721 14223 28779 14229
rect 30282 14220 30288 14232
rect 30340 14220 30346 14272
rect 31846 14260 31852 14272
rect 31807 14232 31852 14260
rect 31846 14220 31852 14232
rect 31904 14220 31910 14272
rect 33410 14260 33416 14272
rect 33371 14232 33416 14260
rect 33410 14220 33416 14232
rect 33468 14220 33474 14272
rect 34606 14220 34612 14272
rect 34664 14260 34670 14272
rect 35621 14263 35679 14269
rect 35621 14260 35633 14263
rect 34664 14232 35633 14260
rect 34664 14220 34670 14232
rect 35621 14229 35633 14232
rect 35667 14260 35679 14263
rect 35866 14260 35894 14436
rect 36262 14424 36268 14436
rect 36320 14424 36326 14476
rect 36449 14467 36507 14473
rect 36449 14433 36461 14467
rect 36495 14464 36507 14467
rect 36538 14464 36544 14476
rect 36495 14436 36544 14464
rect 36495 14433 36507 14436
rect 36449 14427 36507 14433
rect 36538 14424 36544 14436
rect 36596 14424 36602 14476
rect 35667 14232 35894 14260
rect 35667 14229 35679 14232
rect 35621 14223 35679 14229
rect 36538 14220 36544 14272
rect 36596 14260 36602 14272
rect 36909 14263 36967 14269
rect 36596 14232 36641 14260
rect 36596 14220 36602 14232
rect 36909 14229 36921 14263
rect 36955 14260 36967 14263
rect 37274 14260 37280 14272
rect 36955 14232 37280 14260
rect 36955 14229 36967 14232
rect 36909 14223 36967 14229
rect 37274 14220 37280 14232
rect 37332 14220 37338 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 16853 14059 16911 14065
rect 16853 14025 16865 14059
rect 16899 14056 16911 14059
rect 17034 14056 17040 14068
rect 16899 14028 17040 14056
rect 16899 14025 16911 14028
rect 16853 14019 16911 14025
rect 17034 14016 17040 14028
rect 17092 14016 17098 14068
rect 18138 14016 18144 14068
rect 18196 14056 18202 14068
rect 18690 14056 18696 14068
rect 18196 14028 18696 14056
rect 18196 14016 18202 14028
rect 18690 14016 18696 14028
rect 18748 14056 18754 14068
rect 23750 14056 23756 14068
rect 18748 14028 23756 14056
rect 18748 14016 18754 14028
rect 23750 14016 23756 14028
rect 23808 14016 23814 14068
rect 25406 14056 25412 14068
rect 25367 14028 25412 14056
rect 25406 14016 25412 14028
rect 25464 14016 25470 14068
rect 25498 14016 25504 14068
rect 25556 14056 25562 14068
rect 31846 14056 31852 14068
rect 25556 14028 31852 14056
rect 25556 14016 25562 14028
rect 31846 14016 31852 14028
rect 31904 14016 31910 14068
rect 20990 13948 20996 14000
rect 21048 13988 21054 14000
rect 27430 13988 27436 14000
rect 21048 13960 27436 13988
rect 21048 13948 21054 13960
rect 27430 13948 27436 13960
rect 27488 13948 27494 14000
rect 15654 13880 15660 13932
rect 15712 13920 15718 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 15712 13892 16681 13920
rect 15712 13880 15718 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 17681 13923 17739 13929
rect 17681 13889 17693 13923
rect 17727 13920 17739 13923
rect 18506 13920 18512 13932
rect 17727 13892 18512 13920
rect 17727 13889 17739 13892
rect 17681 13883 17739 13889
rect 18506 13880 18512 13892
rect 18564 13880 18570 13932
rect 20162 13920 20168 13932
rect 20123 13892 20168 13920
rect 20162 13880 20168 13892
rect 20220 13880 20226 13932
rect 20349 13923 20407 13929
rect 20349 13889 20361 13923
rect 20395 13920 20407 13923
rect 21082 13920 21088 13932
rect 20395 13892 21088 13920
rect 20395 13889 20407 13892
rect 20349 13883 20407 13889
rect 21082 13880 21088 13892
rect 21140 13920 21146 13932
rect 22646 13920 22652 13932
rect 21140 13892 22652 13920
rect 21140 13880 21146 13892
rect 22646 13880 22652 13892
rect 22704 13880 22710 13932
rect 25406 13880 25412 13932
rect 25464 13920 25470 13932
rect 30098 13920 30104 13932
rect 25464 13892 30104 13920
rect 25464 13880 25470 13892
rect 30098 13880 30104 13892
rect 30156 13880 30162 13932
rect 36446 13920 36452 13932
rect 36407 13892 36452 13920
rect 36446 13880 36452 13892
rect 36504 13880 36510 13932
rect 15838 13852 15844 13864
rect 15751 13824 15844 13852
rect 15838 13812 15844 13824
rect 15896 13852 15902 13864
rect 17402 13852 17408 13864
rect 15896 13824 17408 13852
rect 15896 13812 15902 13824
rect 17402 13812 17408 13824
rect 17460 13852 17466 13864
rect 17497 13855 17555 13861
rect 17497 13852 17509 13855
rect 17460 13824 17509 13852
rect 17460 13812 17466 13824
rect 17497 13821 17509 13824
rect 17543 13821 17555 13855
rect 17497 13815 17555 13821
rect 17865 13855 17923 13861
rect 17865 13821 17877 13855
rect 17911 13852 17923 13855
rect 18230 13852 18236 13864
rect 17911 13824 18236 13852
rect 17911 13821 17923 13824
rect 17865 13815 17923 13821
rect 18230 13812 18236 13824
rect 18288 13812 18294 13864
rect 20254 13812 20260 13864
rect 20312 13852 20318 13864
rect 25498 13852 25504 13864
rect 20312 13824 25504 13852
rect 20312 13812 20318 13824
rect 25498 13812 25504 13824
rect 25556 13812 25562 13864
rect 20990 13744 20996 13796
rect 21048 13784 21054 13796
rect 22186 13784 22192 13796
rect 21048 13756 22192 13784
rect 21048 13744 21054 13756
rect 22186 13744 22192 13756
rect 22244 13744 22250 13796
rect 23750 13744 23756 13796
rect 23808 13784 23814 13796
rect 30374 13784 30380 13796
rect 23808 13756 30380 13784
rect 23808 13744 23814 13756
rect 30374 13744 30380 13756
rect 30432 13744 30438 13796
rect 19886 13676 19892 13728
rect 19944 13716 19950 13728
rect 19981 13719 20039 13725
rect 19981 13716 19993 13719
rect 19944 13688 19993 13716
rect 19944 13676 19950 13688
rect 19981 13685 19993 13688
rect 20027 13685 20039 13719
rect 36262 13716 36268 13728
rect 36223 13688 36268 13716
rect 19981 13679 20039 13685
rect 36262 13676 36268 13688
rect 36320 13676 36326 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 19429 13515 19487 13521
rect 19429 13481 19441 13515
rect 19475 13512 19487 13515
rect 19475 13484 26234 13512
rect 19475 13481 19487 13484
rect 19429 13475 19487 13481
rect 18046 13404 18052 13456
rect 18104 13444 18110 13456
rect 21637 13447 21695 13453
rect 21637 13444 21649 13447
rect 18104 13416 21649 13444
rect 18104 13404 18110 13416
rect 21637 13413 21649 13416
rect 21683 13413 21695 13447
rect 24486 13444 24492 13456
rect 24447 13416 24492 13444
rect 21637 13407 21695 13413
rect 24486 13404 24492 13416
rect 24544 13404 24550 13456
rect 14366 13308 14372 13320
rect 14327 13280 14372 13308
rect 14366 13268 14372 13280
rect 14424 13268 14430 13320
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13308 15623 13311
rect 16117 13311 16175 13317
rect 16117 13308 16129 13311
rect 15611 13280 16129 13308
rect 15611 13277 15623 13280
rect 15565 13271 15623 13277
rect 16117 13277 16129 13280
rect 16163 13308 16175 13311
rect 16666 13308 16672 13320
rect 16163 13280 16672 13308
rect 16163 13277 16175 13280
rect 16117 13271 16175 13277
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 16761 13311 16819 13317
rect 16761 13277 16773 13311
rect 16807 13308 16819 13311
rect 17770 13308 17776 13320
rect 16807 13280 17776 13308
rect 16807 13277 16819 13280
rect 16761 13271 16819 13277
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 18230 13308 18236 13320
rect 18191 13280 18236 13308
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 19242 13308 19248 13320
rect 19203 13280 19248 13308
rect 19242 13268 19248 13280
rect 19300 13268 19306 13320
rect 19886 13308 19892 13320
rect 19847 13280 19892 13308
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 23014 13308 23020 13320
rect 22975 13280 23020 13308
rect 23014 13268 23020 13280
rect 23072 13268 23078 13320
rect 25866 13308 25872 13320
rect 25827 13280 25872 13308
rect 25866 13268 25872 13280
rect 25924 13268 25930 13320
rect 22750 13243 22808 13249
rect 22750 13240 22762 13243
rect 18248 13212 22762 13240
rect 18248 13184 18276 13212
rect 22750 13209 22762 13212
rect 22796 13209 22808 13243
rect 22750 13203 22808 13209
rect 22922 13200 22928 13252
rect 22980 13240 22986 13252
rect 25602 13243 25660 13249
rect 25602 13240 25614 13243
rect 22980 13212 25614 13240
rect 22980 13200 22986 13212
rect 25602 13209 25614 13212
rect 25648 13209 25660 13243
rect 26206 13240 26234 13484
rect 36630 13472 36636 13524
rect 36688 13512 36694 13524
rect 36725 13515 36783 13521
rect 36725 13512 36737 13515
rect 36688 13484 36737 13512
rect 36688 13472 36694 13484
rect 36725 13481 36737 13484
rect 36771 13481 36783 13515
rect 36725 13475 36783 13481
rect 27154 13268 27160 13320
rect 27212 13308 27218 13320
rect 27709 13311 27767 13317
rect 27709 13308 27721 13311
rect 27212 13280 27721 13308
rect 27212 13268 27218 13280
rect 27709 13277 27721 13280
rect 27755 13277 27767 13311
rect 27709 13271 27767 13277
rect 31754 13268 31760 13320
rect 31812 13308 31818 13320
rect 32585 13311 32643 13317
rect 32585 13308 32597 13311
rect 31812 13280 32597 13308
rect 31812 13268 31818 13280
rect 32585 13277 32597 13280
rect 32631 13277 32643 13311
rect 38102 13308 38108 13320
rect 38063 13280 38108 13308
rect 32585 13271 32643 13277
rect 38102 13268 38108 13280
rect 38160 13268 38166 13320
rect 27442 13243 27500 13249
rect 27442 13240 27454 13243
rect 26206 13212 27454 13240
rect 25602 13203 25660 13209
rect 27442 13209 27454 13212
rect 27488 13209 27500 13243
rect 27442 13203 27500 13209
rect 30282 13200 30288 13252
rect 30340 13240 30346 13252
rect 32318 13243 32376 13249
rect 32318 13240 32330 13243
rect 30340 13212 32330 13240
rect 30340 13200 30346 13212
rect 32318 13209 32330 13212
rect 32364 13209 32376 13243
rect 32318 13203 32376 13209
rect 37458 13200 37464 13252
rect 37516 13240 37522 13252
rect 37838 13243 37896 13249
rect 37838 13240 37850 13243
rect 37516 13212 37850 13240
rect 37516 13200 37522 13212
rect 37838 13209 37850 13212
rect 37884 13209 37896 13243
rect 37838 13203 37896 13209
rect 14550 13172 14556 13184
rect 14511 13144 14556 13172
rect 14550 13132 14556 13144
rect 14608 13132 14614 13184
rect 16945 13175 17003 13181
rect 16945 13141 16957 13175
rect 16991 13172 17003 13175
rect 17310 13172 17316 13184
rect 16991 13144 17316 13172
rect 16991 13141 17003 13144
rect 16945 13135 17003 13141
rect 17310 13132 17316 13144
rect 17368 13132 17374 13184
rect 17402 13132 17408 13184
rect 17460 13172 17466 13184
rect 17497 13175 17555 13181
rect 17497 13172 17509 13175
rect 17460 13144 17509 13172
rect 17460 13132 17466 13144
rect 17497 13141 17509 13144
rect 17543 13172 17555 13175
rect 17770 13172 17776 13184
rect 17543 13144 17776 13172
rect 17543 13141 17555 13144
rect 17497 13135 17555 13141
rect 17770 13132 17776 13144
rect 17828 13132 17834 13184
rect 18230 13132 18236 13184
rect 18288 13132 18294 13184
rect 18414 13172 18420 13184
rect 18375 13144 18420 13172
rect 18414 13132 18420 13144
rect 18472 13132 18478 13184
rect 20070 13172 20076 13184
rect 20031 13144 20076 13172
rect 20070 13132 20076 13144
rect 20128 13132 20134 13184
rect 22186 13132 22192 13184
rect 22244 13172 22250 13184
rect 26329 13175 26387 13181
rect 26329 13172 26341 13175
rect 22244 13144 26341 13172
rect 22244 13132 22250 13144
rect 26329 13141 26341 13144
rect 26375 13141 26387 13175
rect 26329 13135 26387 13141
rect 30098 13132 30104 13184
rect 30156 13172 30162 13184
rect 31205 13175 31263 13181
rect 31205 13172 31217 13175
rect 30156 13144 31217 13172
rect 30156 13132 30162 13144
rect 31205 13141 31217 13144
rect 31251 13141 31263 13175
rect 31205 13135 31263 13141
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 14550 12928 14556 12980
rect 14608 12968 14614 12980
rect 22922 12968 22928 12980
rect 14608 12940 22928 12968
rect 14608 12928 14614 12940
rect 22922 12928 22928 12940
rect 22980 12928 22986 12980
rect 32122 12968 32128 12980
rect 32083 12940 32128 12968
rect 32122 12928 32128 12940
rect 32180 12928 32186 12980
rect 33778 12928 33784 12980
rect 33836 12968 33842 12980
rect 33965 12971 34023 12977
rect 33965 12968 33977 12971
rect 33836 12940 33977 12968
rect 33836 12928 33842 12940
rect 33965 12937 33977 12940
rect 34011 12937 34023 12971
rect 37458 12968 37464 12980
rect 37419 12940 37464 12968
rect 33965 12931 34023 12937
rect 37458 12928 37464 12940
rect 37516 12928 37522 12980
rect 16117 12903 16175 12909
rect 16117 12869 16129 12903
rect 16163 12900 16175 12903
rect 16163 12872 17540 12900
rect 16163 12869 16175 12872
rect 16117 12863 16175 12869
rect 15930 12832 15936 12844
rect 15891 12804 15936 12832
rect 15930 12792 15936 12804
rect 15988 12792 15994 12844
rect 16850 12832 16856 12844
rect 16811 12804 16856 12832
rect 16850 12792 16856 12804
rect 16908 12792 16914 12844
rect 17512 12841 17540 12872
rect 18414 12860 18420 12912
rect 18472 12900 18478 12912
rect 18472 12872 26234 12900
rect 18472 12860 18478 12872
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12801 17555 12835
rect 18966 12832 18972 12844
rect 18927 12804 18972 12832
rect 17497 12795 17555 12801
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 19797 12835 19855 12841
rect 19797 12801 19809 12835
rect 19843 12832 19855 12835
rect 19978 12832 19984 12844
rect 19843 12804 19984 12832
rect 19843 12801 19855 12804
rect 19797 12795 19855 12801
rect 19978 12792 19984 12804
rect 20036 12792 20042 12844
rect 20625 12835 20683 12841
rect 20625 12801 20637 12835
rect 20671 12832 20683 12835
rect 20714 12832 20720 12844
rect 20671 12804 20720 12832
rect 20671 12801 20683 12804
rect 20625 12795 20683 12801
rect 20714 12792 20720 12804
rect 20772 12792 20778 12844
rect 20898 12792 20904 12844
rect 20956 12832 20962 12844
rect 22934 12835 22992 12841
rect 22934 12832 22946 12835
rect 20956 12804 22946 12832
rect 20956 12792 20962 12804
rect 22934 12801 22946 12804
rect 22980 12801 22992 12835
rect 22934 12795 22992 12801
rect 23750 12792 23756 12844
rect 23808 12832 23814 12844
rect 24774 12835 24832 12841
rect 24774 12832 24786 12835
rect 23808 12804 24786 12832
rect 23808 12792 23814 12804
rect 24774 12801 24786 12804
rect 24820 12801 24832 12835
rect 24774 12795 24832 12801
rect 25041 12835 25099 12841
rect 25041 12801 25053 12835
rect 25087 12832 25099 12835
rect 25498 12832 25504 12844
rect 25087 12804 25504 12832
rect 25087 12801 25099 12804
rect 25041 12795 25099 12801
rect 25498 12792 25504 12804
rect 25556 12832 25562 12844
rect 25866 12832 25872 12844
rect 25556 12804 25872 12832
rect 25556 12792 25562 12804
rect 25866 12792 25872 12804
rect 25924 12792 25930 12844
rect 26206 12832 26234 12872
rect 27154 12860 27160 12912
rect 27212 12900 27218 12912
rect 27212 12872 28948 12900
rect 27212 12860 27218 12872
rect 28920 12841 28948 12872
rect 29546 12860 29552 12912
rect 29604 12900 29610 12912
rect 30478 12903 30536 12909
rect 30478 12900 30490 12903
rect 29604 12872 30490 12900
rect 29604 12860 29610 12872
rect 30478 12869 30490 12872
rect 30524 12869 30536 12903
rect 30478 12863 30536 12869
rect 33260 12903 33318 12909
rect 33260 12869 33272 12903
rect 33306 12900 33318 12903
rect 33410 12900 33416 12912
rect 33306 12872 33416 12900
rect 33306 12869 33318 12872
rect 33260 12863 33318 12869
rect 33410 12860 33416 12872
rect 33468 12860 33474 12912
rect 33520 12872 35388 12900
rect 33520 12841 33548 12872
rect 35360 12844 35388 12872
rect 28638 12835 28696 12841
rect 28638 12832 28650 12835
rect 26206 12804 28650 12832
rect 28638 12801 28650 12804
rect 28684 12801 28696 12835
rect 28638 12795 28696 12801
rect 28905 12835 28963 12841
rect 28905 12801 28917 12835
rect 28951 12801 28963 12835
rect 28905 12795 28963 12801
rect 33505 12835 33563 12841
rect 33505 12801 33517 12835
rect 33551 12801 33563 12835
rect 33505 12795 33563 12801
rect 34790 12792 34796 12844
rect 34848 12832 34854 12844
rect 35078 12835 35136 12841
rect 35078 12832 35090 12835
rect 34848 12804 35090 12832
rect 34848 12792 34854 12804
rect 35078 12801 35090 12804
rect 35124 12801 35136 12835
rect 35342 12832 35348 12844
rect 35255 12804 35348 12832
rect 35078 12795 35136 12801
rect 35342 12792 35348 12804
rect 35400 12792 35406 12844
rect 37274 12832 37280 12844
rect 37235 12804 37280 12832
rect 37274 12792 37280 12804
rect 37332 12792 37338 12844
rect 15289 12767 15347 12773
rect 15289 12733 15301 12767
rect 15335 12764 15347 12767
rect 15749 12767 15807 12773
rect 15749 12764 15761 12767
rect 15335 12736 15761 12764
rect 15335 12733 15347 12736
rect 15289 12727 15347 12733
rect 15749 12733 15761 12736
rect 15795 12764 15807 12767
rect 16666 12764 16672 12776
rect 15795 12736 16672 12764
rect 15795 12733 15807 12736
rect 15749 12727 15807 12733
rect 16666 12724 16672 12736
rect 16724 12764 16730 12776
rect 17770 12764 17776 12776
rect 16724 12736 17776 12764
rect 16724 12724 16730 12736
rect 17770 12724 17776 12736
rect 17828 12764 17834 12776
rect 18325 12767 18383 12773
rect 18325 12764 18337 12767
rect 17828 12736 18337 12764
rect 17828 12724 17834 12736
rect 18325 12733 18337 12736
rect 18371 12764 18383 12767
rect 18782 12764 18788 12776
rect 18371 12736 18788 12764
rect 18371 12733 18383 12736
rect 18325 12727 18383 12733
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12764 19671 12767
rect 19886 12764 19892 12776
rect 19659 12736 19892 12764
rect 19659 12733 19671 12736
rect 19613 12727 19671 12733
rect 19886 12724 19892 12736
rect 19944 12764 19950 12776
rect 20809 12767 20867 12773
rect 20809 12764 20821 12767
rect 19944 12736 20821 12764
rect 19944 12724 19950 12736
rect 20809 12733 20821 12736
rect 20855 12764 20867 12767
rect 21082 12764 21088 12776
rect 20855 12736 21088 12764
rect 20855 12733 20867 12736
rect 20809 12727 20867 12733
rect 21082 12724 21088 12736
rect 21140 12724 21146 12776
rect 21174 12724 21180 12776
rect 21232 12764 21238 12776
rect 21818 12764 21824 12776
rect 21232 12736 21824 12764
rect 21232 12724 21238 12736
rect 21818 12724 21824 12736
rect 21876 12764 21882 12776
rect 23198 12764 23204 12776
rect 21876 12736 22094 12764
rect 23159 12736 23204 12764
rect 21876 12724 21882 12736
rect 17681 12699 17739 12705
rect 17681 12665 17693 12699
rect 17727 12696 17739 12699
rect 20622 12696 20628 12708
rect 17727 12668 20628 12696
rect 17727 12665 17739 12668
rect 17681 12659 17739 12665
rect 20622 12656 20628 12668
rect 20680 12656 20686 12708
rect 22066 12696 22094 12736
rect 23198 12724 23204 12736
rect 23256 12724 23262 12776
rect 30745 12767 30803 12773
rect 30745 12733 30757 12767
rect 30791 12764 30803 12767
rect 31754 12764 31760 12776
rect 30791 12736 31760 12764
rect 30791 12733 30803 12736
rect 30745 12727 30803 12733
rect 31754 12724 31760 12736
rect 31812 12724 31818 12776
rect 22066 12668 22324 12696
rect 17037 12631 17095 12637
rect 17037 12597 17049 12631
rect 17083 12628 17095 12631
rect 17218 12628 17224 12640
rect 17083 12600 17224 12628
rect 17083 12597 17095 12600
rect 17037 12591 17095 12597
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 19153 12631 19211 12637
rect 19153 12597 19165 12631
rect 19199 12628 19211 12631
rect 19242 12628 19248 12640
rect 19199 12600 19248 12628
rect 19199 12597 19211 12600
rect 19153 12591 19211 12597
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 19981 12631 20039 12637
rect 19981 12597 19993 12631
rect 20027 12628 20039 12631
rect 20070 12628 20076 12640
rect 20027 12600 20076 12628
rect 20027 12597 20039 12600
rect 19981 12591 20039 12597
rect 20070 12588 20076 12600
rect 20128 12588 20134 12640
rect 20438 12628 20444 12640
rect 20399 12600 20444 12628
rect 20438 12588 20444 12600
rect 20496 12588 20502 12640
rect 21818 12628 21824 12640
rect 21779 12600 21824 12628
rect 21818 12588 21824 12600
rect 21876 12588 21882 12640
rect 22296 12628 22324 12668
rect 23492 12668 23796 12696
rect 23492 12628 23520 12668
rect 23658 12628 23664 12640
rect 22296 12600 23520 12628
rect 23619 12600 23664 12628
rect 23658 12588 23664 12600
rect 23716 12588 23722 12640
rect 23768 12628 23796 12668
rect 27246 12656 27252 12708
rect 27304 12696 27310 12708
rect 27304 12668 27844 12696
rect 27304 12656 27310 12668
rect 27525 12631 27583 12637
rect 27525 12628 27537 12631
rect 23768 12600 27537 12628
rect 27525 12597 27537 12600
rect 27571 12597 27583 12631
rect 27816 12628 27844 12668
rect 29365 12631 29423 12637
rect 29365 12628 29377 12631
rect 27816 12600 29377 12628
rect 27525 12591 27583 12597
rect 29365 12597 29377 12600
rect 29411 12597 29423 12631
rect 29365 12591 29423 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 13170 12384 13176 12436
rect 13228 12424 13234 12436
rect 13722 12424 13728 12436
rect 13228 12396 13728 12424
rect 13228 12384 13234 12396
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 18230 12384 18236 12436
rect 18288 12424 18294 12436
rect 18325 12427 18383 12433
rect 18325 12424 18337 12427
rect 18288 12396 18337 12424
rect 18288 12384 18294 12396
rect 18325 12393 18337 12396
rect 18371 12393 18383 12427
rect 18325 12387 18383 12393
rect 18782 12384 18788 12436
rect 18840 12424 18846 12436
rect 20073 12427 20131 12433
rect 20073 12424 20085 12427
rect 18840 12396 20085 12424
rect 18840 12384 18846 12396
rect 20073 12393 20085 12396
rect 20119 12424 20131 12427
rect 20254 12424 20260 12436
rect 20119 12396 20260 12424
rect 20119 12393 20131 12396
rect 20073 12387 20131 12393
rect 20254 12384 20260 12396
rect 20312 12384 20318 12436
rect 21634 12424 21640 12436
rect 21595 12396 21640 12424
rect 21634 12384 21640 12396
rect 21692 12384 21698 12436
rect 25777 12427 25835 12433
rect 25777 12424 25789 12427
rect 22066 12396 25789 12424
rect 17494 12316 17500 12368
rect 17552 12356 17558 12368
rect 17770 12356 17776 12368
rect 17552 12328 17776 12356
rect 17552 12316 17558 12328
rect 17770 12316 17776 12328
rect 17828 12356 17834 12368
rect 22066 12356 22094 12396
rect 25777 12393 25789 12396
rect 25823 12393 25835 12427
rect 25777 12387 25835 12393
rect 37366 12384 37372 12436
rect 37424 12424 37430 12436
rect 37461 12427 37519 12433
rect 37461 12424 37473 12427
rect 37424 12396 37473 12424
rect 37424 12384 37430 12396
rect 37461 12393 37473 12396
rect 37507 12393 37519 12427
rect 37461 12387 37519 12393
rect 17828 12328 22094 12356
rect 17828 12316 17834 12328
rect 15473 12291 15531 12297
rect 15473 12257 15485 12291
rect 15519 12288 15531 12291
rect 15519 12260 16896 12288
rect 15519 12257 15531 12260
rect 15473 12251 15531 12257
rect 14921 12223 14979 12229
rect 14921 12189 14933 12223
rect 14967 12220 14979 12223
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 14967 12192 15945 12220
rect 14967 12189 14979 12192
rect 14921 12183 14979 12189
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 16117 12223 16175 12229
rect 16117 12189 16129 12223
rect 16163 12220 16175 12223
rect 16574 12220 16580 12232
rect 16163 12192 16580 12220
rect 16163 12189 16175 12192
rect 16117 12183 16175 12189
rect 15948 12152 15976 12183
rect 16574 12180 16580 12192
rect 16632 12180 16638 12232
rect 16868 12164 16896 12260
rect 17954 12248 17960 12300
rect 18012 12288 18018 12300
rect 19613 12291 19671 12297
rect 18012 12260 19564 12288
rect 18012 12248 18018 12260
rect 17494 12220 17500 12232
rect 17455 12192 17500 12220
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 18138 12220 18144 12232
rect 18099 12192 18144 12220
rect 18138 12180 18144 12192
rect 18196 12180 18202 12232
rect 19334 12180 19340 12232
rect 19392 12220 19398 12232
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 19392 12192 19441 12220
rect 19392 12180 19398 12192
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 19536 12220 19564 12260
rect 19613 12257 19625 12291
rect 19659 12288 19671 12291
rect 20254 12288 20260 12300
rect 19659 12260 20260 12288
rect 19659 12257 19671 12260
rect 19613 12251 19671 12257
rect 20254 12248 20260 12260
rect 20312 12248 20318 12300
rect 27154 12288 27160 12300
rect 27115 12260 27160 12288
rect 27154 12248 27160 12260
rect 27212 12248 27218 12300
rect 22750 12223 22808 12229
rect 22750 12220 22762 12223
rect 19536 12192 22762 12220
rect 19429 12183 19487 12189
rect 22750 12189 22762 12192
rect 22796 12189 22808 12223
rect 23014 12220 23020 12232
rect 22927 12192 23020 12220
rect 22750 12183 22808 12189
rect 23014 12180 23020 12192
rect 23072 12220 23078 12232
rect 23198 12220 23204 12232
rect 23072 12192 23204 12220
rect 23072 12180 23078 12192
rect 23198 12180 23204 12192
rect 23256 12180 23262 12232
rect 26602 12180 26608 12232
rect 26660 12220 26666 12232
rect 26890 12223 26948 12229
rect 26890 12220 26902 12223
rect 26660 12192 26902 12220
rect 26660 12180 26666 12192
rect 26890 12189 26902 12192
rect 26936 12189 26948 12223
rect 27172 12220 27200 12248
rect 28997 12223 29055 12229
rect 28997 12220 29009 12223
rect 27172 12192 29009 12220
rect 26890 12183 26948 12189
rect 28997 12189 29009 12192
rect 29043 12189 29055 12223
rect 28997 12183 29055 12189
rect 30466 12180 30472 12232
rect 30524 12220 30530 12232
rect 30846 12223 30904 12229
rect 30846 12220 30858 12223
rect 30524 12192 30858 12220
rect 30524 12180 30530 12192
rect 30846 12189 30858 12192
rect 30892 12189 30904 12223
rect 30846 12183 30904 12189
rect 31113 12223 31171 12229
rect 31113 12189 31125 12223
rect 31159 12220 31171 12223
rect 31754 12220 31760 12232
rect 31159 12192 31760 12220
rect 31159 12189 31171 12192
rect 31113 12183 31171 12189
rect 31754 12180 31760 12192
rect 31812 12220 31818 12232
rect 31938 12220 31944 12232
rect 31812 12192 31944 12220
rect 31812 12180 31818 12192
rect 31938 12180 31944 12192
rect 31996 12180 32002 12232
rect 35342 12180 35348 12232
rect 35400 12220 35406 12232
rect 36081 12223 36139 12229
rect 36081 12220 36093 12223
rect 35400 12192 36093 12220
rect 35400 12180 35406 12192
rect 36081 12189 36093 12192
rect 36127 12220 36139 12223
rect 38102 12220 38108 12232
rect 36127 12192 38108 12220
rect 36127 12189 36139 12192
rect 36081 12183 36139 12189
rect 38102 12180 38108 12192
rect 38160 12180 38166 12232
rect 16666 12152 16672 12164
rect 15948 12124 16672 12152
rect 16666 12112 16672 12124
rect 16724 12152 16730 12164
rect 16761 12155 16819 12161
rect 16761 12152 16773 12155
rect 16724 12124 16773 12152
rect 16724 12112 16730 12124
rect 16761 12121 16773 12124
rect 16807 12121 16819 12155
rect 16761 12115 16819 12121
rect 16850 12112 16856 12164
rect 16908 12152 16914 12164
rect 16945 12155 17003 12161
rect 16945 12152 16957 12155
rect 16908 12124 16957 12152
rect 16908 12112 16914 12124
rect 16945 12121 16957 12124
rect 16991 12121 17003 12155
rect 25222 12152 25228 12164
rect 16945 12115 17003 12121
rect 17696 12124 25228 12152
rect 16301 12087 16359 12093
rect 16301 12053 16313 12087
rect 16347 12084 16359 12087
rect 16574 12084 16580 12096
rect 16347 12056 16580 12084
rect 16347 12053 16359 12056
rect 16301 12047 16359 12053
rect 16574 12044 16580 12056
rect 16632 12044 16638 12096
rect 17696 12093 17724 12124
rect 25222 12112 25228 12124
rect 25280 12112 25286 12164
rect 27706 12112 27712 12164
rect 27764 12152 27770 12164
rect 36354 12161 36360 12164
rect 28730 12155 28788 12161
rect 28730 12152 28742 12155
rect 27764 12124 28742 12152
rect 27764 12112 27770 12124
rect 28730 12121 28742 12124
rect 28776 12121 28788 12155
rect 28730 12115 28788 12121
rect 36348 12115 36360 12161
rect 36412 12152 36418 12164
rect 36412 12124 36448 12152
rect 36354 12112 36360 12115
rect 36412 12112 36418 12124
rect 17681 12087 17739 12093
rect 17681 12053 17693 12087
rect 17727 12053 17739 12087
rect 17681 12047 17739 12053
rect 18506 12044 18512 12096
rect 18564 12084 18570 12096
rect 19245 12087 19303 12093
rect 19245 12084 19257 12087
rect 18564 12056 19257 12084
rect 18564 12044 18570 12056
rect 19245 12053 19257 12056
rect 19291 12053 19303 12087
rect 19245 12047 19303 12053
rect 19334 12044 19340 12096
rect 19392 12084 19398 12096
rect 19518 12084 19524 12096
rect 19392 12056 19524 12084
rect 19392 12044 19398 12056
rect 19518 12044 19524 12056
rect 19576 12044 19582 12096
rect 23382 12044 23388 12096
rect 23440 12084 23446 12096
rect 27617 12087 27675 12093
rect 27617 12084 27629 12087
rect 23440 12056 27629 12084
rect 23440 12044 23446 12056
rect 27617 12053 27629 12056
rect 27663 12053 27675 12087
rect 29730 12084 29736 12096
rect 29691 12056 29736 12084
rect 27617 12047 27675 12053
rect 29730 12044 29736 12056
rect 29788 12044 29794 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 17497 11883 17555 11889
rect 17497 11849 17509 11883
rect 17543 11880 17555 11883
rect 18138 11880 18144 11892
rect 17543 11852 18144 11880
rect 17543 11849 17555 11852
rect 17497 11843 17555 11849
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 18601 11883 18659 11889
rect 18601 11849 18613 11883
rect 18647 11880 18659 11883
rect 21450 11880 21456 11892
rect 18647 11852 21456 11880
rect 18647 11849 18659 11852
rect 18601 11843 18659 11849
rect 21450 11840 21456 11852
rect 21508 11880 21514 11892
rect 24121 11883 24179 11889
rect 24121 11880 24133 11883
rect 21508 11852 24133 11880
rect 21508 11840 21514 11852
rect 24121 11849 24133 11852
rect 24167 11849 24179 11883
rect 24121 11843 24179 11849
rect 24228 11852 25452 11880
rect 17037 11815 17095 11821
rect 17037 11781 17049 11815
rect 17083 11812 17095 11815
rect 18046 11812 18052 11824
rect 17083 11784 18052 11812
rect 17083 11781 17095 11784
rect 17037 11775 17095 11781
rect 18046 11772 18052 11784
rect 18104 11812 18110 11824
rect 20165 11815 20223 11821
rect 20165 11812 20177 11815
rect 18104 11784 20177 11812
rect 18104 11772 18110 11784
rect 20165 11781 20177 11784
rect 20211 11781 20223 11815
rect 24228 11812 24256 11852
rect 20165 11775 20223 11781
rect 22066 11784 24256 11812
rect 15562 11744 15568 11756
rect 15523 11716 15568 11744
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 17126 11744 17132 11756
rect 17087 11716 17132 11744
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 18230 11744 18236 11756
rect 17236 11716 18236 11744
rect 15378 11636 15384 11688
rect 15436 11676 15442 11688
rect 16945 11679 17003 11685
rect 16945 11676 16957 11679
rect 15436 11648 16957 11676
rect 15436 11636 15442 11648
rect 16945 11645 16957 11648
rect 16991 11676 17003 11679
rect 17236 11676 17264 11716
rect 18230 11704 18236 11716
rect 18288 11704 18294 11756
rect 18509 11747 18567 11753
rect 18509 11713 18521 11747
rect 18555 11713 18567 11747
rect 18509 11707 18567 11713
rect 19521 11747 19579 11753
rect 19521 11713 19533 11747
rect 19567 11744 19579 11747
rect 20438 11744 20444 11756
rect 19567 11716 20444 11744
rect 19567 11713 19579 11716
rect 19521 11707 19579 11713
rect 16991 11648 17264 11676
rect 16991 11645 17003 11648
rect 16945 11639 17003 11645
rect 18046 11636 18052 11688
rect 18104 11676 18110 11688
rect 18524 11676 18552 11707
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 18104 11648 18552 11676
rect 18693 11679 18751 11685
rect 18104 11636 18110 11648
rect 18693 11645 18705 11679
rect 18739 11645 18751 11679
rect 20898 11676 20904 11688
rect 18693 11639 18751 11645
rect 18800 11648 20904 11676
rect 17494 11568 17500 11620
rect 17552 11608 17558 11620
rect 18141 11611 18199 11617
rect 18141 11608 18153 11611
rect 17552 11580 18153 11608
rect 17552 11568 17558 11580
rect 18141 11577 18153 11580
rect 18187 11577 18199 11611
rect 18141 11571 18199 11577
rect 18230 11568 18236 11620
rect 18288 11608 18294 11620
rect 18708 11608 18736 11639
rect 18288 11580 18736 11608
rect 18288 11568 18294 11580
rect 15749 11543 15807 11549
rect 15749 11509 15761 11543
rect 15795 11540 15807 11543
rect 18800 11540 18828 11648
rect 20898 11636 20904 11648
rect 20956 11636 20962 11688
rect 19334 11568 19340 11620
rect 19392 11608 19398 11620
rect 22066 11608 22094 11784
rect 25222 11772 25228 11824
rect 25280 11821 25286 11824
rect 25280 11812 25292 11821
rect 25424 11812 25452 11852
rect 25590 11840 25596 11892
rect 25648 11880 25654 11892
rect 25648 11852 28580 11880
rect 25648 11840 25654 11852
rect 26326 11812 26332 11824
rect 25280 11784 25325 11812
rect 25424 11784 26332 11812
rect 25280 11775 25292 11784
rect 25280 11772 25286 11775
rect 26326 11772 26332 11784
rect 26384 11772 26390 11824
rect 27154 11772 27160 11824
rect 27212 11812 27218 11824
rect 28552 11812 28580 11852
rect 29178 11840 29184 11892
rect 29236 11880 29242 11892
rect 31754 11880 31760 11892
rect 29236 11852 31760 11880
rect 29236 11840 29242 11852
rect 31754 11840 31760 11852
rect 31812 11880 31818 11892
rect 32217 11883 32275 11889
rect 32217 11880 32229 11883
rect 31812 11852 32229 11880
rect 31812 11840 31818 11852
rect 32217 11849 32229 11852
rect 32263 11849 32275 11883
rect 32217 11843 32275 11849
rect 33330 11815 33388 11821
rect 33330 11812 33342 11815
rect 27212 11784 28488 11812
rect 28552 11784 33342 11812
rect 27212 11772 27218 11784
rect 22186 11704 22192 11756
rect 22244 11744 22250 11756
rect 22934 11747 22992 11753
rect 22934 11744 22946 11747
rect 22244 11716 22946 11744
rect 22244 11704 22250 11716
rect 22934 11713 22946 11716
rect 22980 11713 22992 11747
rect 25498 11744 25504 11756
rect 25459 11716 25504 11744
rect 22934 11707 22992 11713
rect 25498 11704 25504 11716
rect 25556 11704 25562 11756
rect 27614 11704 27620 11756
rect 27672 11744 27678 11756
rect 28460 11753 28488 11784
rect 33330 11781 33342 11784
rect 33376 11781 33388 11815
rect 33330 11775 33388 11781
rect 28178 11747 28236 11753
rect 28178 11744 28190 11747
rect 27672 11716 28190 11744
rect 27672 11704 27678 11716
rect 28178 11713 28190 11716
rect 28224 11713 28236 11747
rect 28178 11707 28236 11713
rect 28445 11747 28503 11753
rect 28445 11713 28457 11747
rect 28491 11713 28503 11747
rect 28445 11707 28503 11713
rect 33597 11747 33655 11753
rect 33597 11713 33609 11747
rect 33643 11744 33655 11747
rect 35342 11744 35348 11756
rect 33643 11716 35348 11744
rect 33643 11713 33655 11716
rect 33597 11707 33655 11713
rect 35342 11704 35348 11716
rect 35400 11704 35406 11756
rect 23198 11676 23204 11688
rect 23159 11648 23204 11676
rect 23198 11636 23204 11648
rect 23256 11636 23262 11688
rect 19392 11580 22094 11608
rect 19392 11568 19398 11580
rect 15795 11512 18828 11540
rect 19705 11543 19763 11549
rect 15795 11509 15807 11512
rect 15749 11503 15807 11509
rect 19705 11509 19717 11543
rect 19751 11540 19763 11543
rect 20438 11540 20444 11552
rect 19751 11512 20444 11540
rect 19751 11509 19763 11512
rect 19705 11503 19763 11509
rect 20438 11500 20444 11512
rect 20496 11500 20502 11552
rect 20530 11500 20536 11552
rect 20588 11540 20594 11552
rect 21821 11543 21879 11549
rect 21821 11540 21833 11543
rect 20588 11512 21833 11540
rect 20588 11500 20594 11512
rect 21821 11509 21833 11512
rect 21867 11540 21879 11543
rect 21910 11540 21916 11552
rect 21867 11512 21916 11540
rect 21867 11509 21879 11512
rect 21821 11503 21879 11509
rect 21910 11500 21916 11512
rect 21968 11500 21974 11552
rect 22462 11500 22468 11552
rect 22520 11540 22526 11552
rect 27065 11543 27123 11549
rect 27065 11540 27077 11543
rect 22520 11512 27077 11540
rect 22520 11500 22526 11512
rect 27065 11509 27077 11512
rect 27111 11509 27123 11543
rect 27065 11503 27123 11509
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 14185 11339 14243 11345
rect 14185 11305 14197 11339
rect 14231 11336 14243 11339
rect 14366 11336 14372 11348
rect 14231 11308 14372 11336
rect 14231 11305 14243 11308
rect 14185 11299 14243 11305
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 14660 11308 15485 11336
rect 13541 11271 13599 11277
rect 13541 11237 13553 11271
rect 13587 11268 13599 11271
rect 13587 11240 14596 11268
rect 13587 11237 13599 11240
rect 13541 11231 13599 11237
rect 13354 11132 13360 11144
rect 13315 11104 13360 11132
rect 13354 11092 13360 11104
rect 13412 11092 13418 11144
rect 14568 11132 14596 11240
rect 14660 11209 14688 11308
rect 15473 11305 15485 11308
rect 15519 11336 15531 11339
rect 16206 11336 16212 11348
rect 15519 11308 16212 11336
rect 15519 11305 15531 11308
rect 15473 11299 15531 11305
rect 16206 11296 16212 11308
rect 16264 11296 16270 11348
rect 17405 11339 17463 11345
rect 17405 11305 17417 11339
rect 17451 11336 17463 11339
rect 17586 11336 17592 11348
rect 17451 11308 17592 11336
rect 17451 11305 17463 11308
rect 17405 11299 17463 11305
rect 17586 11296 17592 11308
rect 17644 11296 17650 11348
rect 18049 11339 18107 11345
rect 18049 11305 18061 11339
rect 18095 11336 18107 11339
rect 30374 11336 30380 11348
rect 18095 11308 27292 11336
rect 30335 11308 30380 11336
rect 18095 11305 18107 11308
rect 18049 11299 18107 11305
rect 16117 11271 16175 11277
rect 16117 11237 16129 11271
rect 16163 11237 16175 11271
rect 16117 11231 16175 11237
rect 16761 11271 16819 11277
rect 16761 11237 16773 11271
rect 16807 11268 16819 11271
rect 17862 11268 17868 11280
rect 16807 11240 17868 11268
rect 16807 11237 16819 11240
rect 16761 11231 16819 11237
rect 14645 11203 14703 11209
rect 14645 11169 14657 11203
rect 14691 11169 14703 11203
rect 14645 11163 14703 11169
rect 14829 11203 14887 11209
rect 14829 11169 14841 11203
rect 14875 11200 14887 11203
rect 15378 11200 15384 11212
rect 14875 11172 15384 11200
rect 14875 11169 14887 11172
rect 14829 11163 14887 11169
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 16132 11200 16160 11231
rect 17862 11228 17868 11240
rect 17920 11228 17926 11280
rect 18693 11271 18751 11277
rect 18693 11237 18705 11271
rect 18739 11268 18751 11271
rect 18739 11240 22094 11268
rect 18739 11237 18751 11240
rect 18693 11231 18751 11237
rect 16132 11172 19656 11200
rect 15194 11132 15200 11144
rect 14568 11104 15200 11132
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 15930 11132 15936 11144
rect 15891 11104 15936 11132
rect 15930 11092 15936 11104
rect 15988 11092 15994 11144
rect 16574 11132 16580 11144
rect 16535 11104 16580 11132
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 17218 11132 17224 11144
rect 17179 11104 17224 11132
rect 17218 11092 17224 11104
rect 17276 11092 17282 11144
rect 17310 11092 17316 11144
rect 17368 11132 17374 11144
rect 17865 11135 17923 11141
rect 17865 11132 17877 11135
rect 17368 11104 17877 11132
rect 17368 11092 17374 11104
rect 17865 11101 17877 11104
rect 17911 11101 17923 11135
rect 18506 11132 18512 11144
rect 18467 11104 18512 11132
rect 17865 11095 17923 11101
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 19242 11132 19248 11144
rect 19203 11104 19248 11132
rect 19242 11092 19248 11104
rect 19300 11092 19306 11144
rect 13630 11024 13636 11076
rect 13688 11064 13694 11076
rect 14553 11067 14611 11073
rect 14553 11064 14565 11067
rect 13688 11036 14565 11064
rect 13688 11024 13694 11036
rect 14553 11033 14565 11036
rect 14599 11033 14611 11067
rect 14553 11027 14611 11033
rect 19334 11024 19340 11076
rect 19392 11064 19398 11076
rect 19628 11064 19656 11172
rect 22066 11132 22094 11240
rect 26605 11203 26663 11209
rect 26605 11169 26617 11203
rect 26651 11200 26663 11203
rect 27154 11200 27160 11212
rect 26651 11172 27160 11200
rect 26651 11169 26663 11172
rect 26605 11163 26663 11169
rect 27154 11160 27160 11172
rect 27212 11160 27218 11212
rect 23109 11135 23167 11141
rect 22066 11104 23060 11132
rect 22842 11067 22900 11073
rect 22842 11064 22854 11067
rect 19392 11036 19472 11064
rect 19628 11036 22854 11064
rect 19392 11024 19398 11036
rect 19444 11005 19472 11036
rect 22842 11033 22854 11036
rect 22888 11033 22900 11067
rect 23032 11064 23060 11104
rect 23109 11101 23121 11135
rect 23155 11132 23167 11135
rect 23198 11132 23204 11144
rect 23155 11104 23204 11132
rect 23155 11101 23167 11104
rect 23109 11095 23167 11101
rect 23198 11092 23204 11104
rect 23256 11092 23262 11144
rect 27264 11132 27292 11308
rect 30374 11296 30380 11308
rect 30432 11296 30438 11348
rect 32582 11296 32588 11348
rect 32640 11336 32646 11348
rect 34701 11339 34759 11345
rect 34701 11336 34713 11339
rect 32640 11308 34713 11336
rect 32640 11296 32646 11308
rect 34701 11305 34713 11308
rect 34747 11305 34759 11339
rect 36725 11339 36783 11345
rect 36725 11336 36737 11339
rect 34701 11299 34759 11305
rect 35084 11308 36737 11336
rect 33318 11228 33324 11280
rect 33376 11268 33382 11280
rect 35084 11268 35112 11308
rect 36725 11305 36737 11308
rect 36771 11305 36783 11339
rect 36725 11299 36783 11305
rect 33376 11240 35112 11268
rect 33376 11228 33382 11240
rect 30006 11160 30012 11212
rect 30064 11200 30070 11212
rect 30742 11200 30748 11212
rect 30064 11172 30748 11200
rect 30064 11160 30070 11172
rect 30742 11160 30748 11172
rect 30800 11160 30806 11212
rect 38102 11200 38108 11212
rect 38063 11172 38108 11200
rect 38102 11160 38108 11172
rect 38160 11160 38166 11212
rect 31490 11135 31548 11141
rect 31490 11132 31502 11135
rect 27264 11104 31502 11132
rect 31490 11101 31502 11104
rect 31536 11101 31548 11135
rect 31490 11095 31548 11101
rect 31757 11135 31815 11141
rect 31757 11101 31769 11135
rect 31803 11132 31815 11135
rect 31938 11132 31944 11144
rect 31803 11104 31944 11132
rect 31803 11101 31815 11104
rect 31757 11095 31815 11101
rect 31938 11092 31944 11104
rect 31996 11132 32002 11144
rect 32217 11135 32275 11141
rect 32217 11132 32229 11135
rect 31996 11104 32229 11132
rect 31996 11092 32002 11104
rect 32217 11101 32229 11104
rect 32263 11101 32275 11135
rect 32217 11095 32275 11101
rect 35526 11092 35532 11144
rect 35584 11132 35590 11144
rect 36081 11135 36139 11141
rect 36081 11132 36093 11135
rect 35584 11104 36093 11132
rect 35584 11092 35590 11104
rect 36081 11101 36093 11104
rect 36127 11132 36139 11135
rect 38120 11132 38148 11160
rect 36127 11104 38148 11132
rect 36127 11101 36139 11104
rect 36081 11095 36139 11101
rect 24762 11064 24768 11076
rect 23032 11036 24768 11064
rect 22842 11027 22900 11033
rect 24762 11024 24768 11036
rect 24820 11024 24826 11076
rect 26234 11024 26240 11076
rect 26292 11064 26298 11076
rect 26338 11067 26396 11073
rect 26338 11064 26350 11067
rect 26292 11036 26350 11064
rect 26292 11024 26298 11036
rect 26338 11033 26350 11036
rect 26384 11033 26396 11067
rect 26338 11027 26396 11033
rect 30650 11024 30656 11076
rect 30708 11064 30714 11076
rect 32462 11067 32520 11073
rect 32462 11064 32474 11067
rect 30708 11036 32474 11064
rect 30708 11024 30714 11036
rect 32462 11033 32474 11036
rect 32508 11033 32520 11067
rect 32462 11027 32520 11033
rect 32674 11024 32680 11076
rect 32732 11064 32738 11076
rect 35814 11067 35872 11073
rect 35814 11064 35826 11067
rect 32732 11036 35826 11064
rect 32732 11024 32738 11036
rect 35814 11033 35826 11036
rect 35860 11033 35872 11067
rect 37826 11064 37832 11076
rect 37884 11073 37890 11076
rect 37796 11036 37832 11064
rect 35814 11027 35872 11033
rect 37826 11024 37832 11036
rect 37884 11027 37896 11073
rect 37884 11024 37890 11027
rect 19429 10999 19487 11005
rect 19429 10965 19441 10999
rect 19475 10965 19487 10999
rect 21726 10996 21732 11008
rect 21687 10968 21732 10996
rect 19429 10959 19487 10965
rect 21726 10956 21732 10968
rect 21784 10956 21790 11008
rect 25222 10996 25228 11008
rect 25183 10968 25228 10996
rect 25222 10956 25228 10968
rect 25280 10956 25286 11008
rect 33597 10999 33655 11005
rect 33597 10965 33609 10999
rect 33643 10996 33655 10999
rect 33686 10996 33692 11008
rect 33643 10968 33692 10996
rect 33643 10965 33655 10968
rect 33597 10959 33655 10965
rect 33686 10956 33692 10968
rect 33744 10996 33750 11008
rect 34238 10996 34244 11008
rect 33744 10968 34244 10996
rect 33744 10956 33750 10968
rect 34238 10956 34244 10968
rect 34296 10956 34302 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 15562 10752 15568 10804
rect 15620 10792 15626 10804
rect 15841 10795 15899 10801
rect 15841 10792 15853 10795
rect 15620 10764 15853 10792
rect 15620 10752 15626 10764
rect 15841 10761 15853 10764
rect 15887 10761 15899 10795
rect 15841 10755 15899 10761
rect 19429 10795 19487 10801
rect 19429 10761 19441 10795
rect 19475 10792 19487 10795
rect 19794 10792 19800 10804
rect 19475 10764 19800 10792
rect 19475 10761 19487 10764
rect 19429 10755 19487 10761
rect 19794 10752 19800 10764
rect 19852 10792 19858 10804
rect 19978 10792 19984 10804
rect 19852 10764 19984 10792
rect 19852 10752 19858 10764
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 30190 10792 30196 10804
rect 21928 10764 30196 10792
rect 15381 10727 15439 10733
rect 15381 10693 15393 10727
rect 15427 10724 15439 10727
rect 15746 10724 15752 10736
rect 15427 10696 15752 10724
rect 15427 10693 15439 10696
rect 15381 10687 15439 10693
rect 15746 10684 15752 10696
rect 15804 10724 15810 10736
rect 16761 10727 16819 10733
rect 16761 10724 16773 10727
rect 15804 10696 16773 10724
rect 15804 10684 15810 10696
rect 16761 10693 16773 10696
rect 16807 10724 16819 10727
rect 21818 10724 21824 10736
rect 16807 10696 21824 10724
rect 16807 10693 16819 10696
rect 16761 10687 16819 10693
rect 21818 10684 21824 10696
rect 21876 10684 21882 10736
rect 11514 10656 11520 10668
rect 11475 10628 11520 10656
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 15470 10656 15476 10668
rect 15431 10628 15476 10656
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10656 18107 10659
rect 18322 10656 18328 10668
rect 18095 10628 18328 10656
rect 18095 10625 18107 10628
rect 18049 10619 18107 10625
rect 18322 10616 18328 10628
rect 18380 10616 18386 10668
rect 19337 10659 19395 10665
rect 19337 10625 19349 10659
rect 19383 10656 19395 10659
rect 20070 10656 20076 10668
rect 19383 10628 19417 10656
rect 20031 10628 20076 10656
rect 19383 10625 19395 10628
rect 19337 10619 19395 10625
rect 15289 10591 15347 10597
rect 15289 10557 15301 10591
rect 15335 10588 15347 10591
rect 15378 10588 15384 10600
rect 15335 10560 15384 10588
rect 15335 10557 15347 10560
rect 15289 10551 15347 10557
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 15562 10548 15568 10600
rect 15620 10588 15626 10600
rect 16850 10588 16856 10600
rect 15620 10560 16856 10588
rect 15620 10548 15626 10560
rect 16850 10548 16856 10560
rect 16908 10588 16914 10600
rect 18785 10591 18843 10597
rect 18785 10588 18797 10591
rect 16908 10560 18797 10588
rect 16908 10548 16914 10560
rect 18785 10557 18797 10560
rect 18831 10588 18843 10591
rect 19352 10588 19380 10619
rect 20070 10616 20076 10628
rect 20128 10616 20134 10668
rect 21928 10588 21956 10764
rect 30190 10752 30196 10764
rect 30248 10752 30254 10804
rect 35526 10724 35532 10736
rect 35487 10696 35532 10724
rect 35526 10684 35532 10696
rect 35584 10684 35590 10736
rect 25133 10659 25191 10665
rect 25133 10625 25145 10659
rect 25179 10656 25191 10659
rect 26050 10656 26056 10668
rect 25179 10628 26056 10656
rect 25179 10625 25191 10628
rect 25133 10619 25191 10625
rect 26050 10616 26056 10628
rect 26108 10616 26114 10668
rect 27154 10616 27160 10668
rect 27212 10656 27218 10668
rect 28350 10656 28356 10668
rect 27212 10628 28356 10656
rect 27212 10616 27218 10628
rect 28350 10616 28356 10628
rect 28408 10656 28414 10668
rect 28537 10659 28595 10665
rect 28537 10656 28549 10659
rect 28408 10628 28549 10656
rect 28408 10616 28414 10628
rect 28537 10625 28549 10628
rect 28583 10625 28595 10659
rect 28793 10659 28851 10665
rect 28793 10656 28805 10659
rect 28537 10619 28595 10625
rect 28644 10628 28805 10656
rect 27614 10588 27620 10600
rect 18831 10560 21956 10588
rect 23124 10560 27620 10588
rect 18831 10557 18843 10560
rect 18785 10551 18843 10557
rect 11698 10520 11704 10532
rect 11659 10492 11704 10520
rect 11698 10480 11704 10492
rect 11756 10480 11762 10532
rect 18233 10523 18291 10529
rect 18233 10489 18245 10523
rect 18279 10520 18291 10523
rect 23124 10520 23152 10560
rect 27614 10548 27620 10560
rect 27672 10548 27678 10600
rect 28644 10588 28672 10628
rect 28793 10625 28805 10628
rect 28839 10625 28851 10659
rect 33778 10656 33784 10668
rect 33739 10628 33784 10656
rect 28793 10619 28851 10625
rect 33778 10616 33784 10628
rect 33836 10616 33842 10668
rect 28552 10560 28672 10588
rect 18279 10492 23152 10520
rect 18279 10489 18291 10492
rect 18233 10483 18291 10489
rect 23198 10480 23204 10532
rect 23256 10520 23262 10532
rect 23845 10523 23903 10529
rect 23845 10520 23857 10523
rect 23256 10492 23857 10520
rect 23256 10480 23262 10492
rect 23845 10489 23857 10492
rect 23891 10520 23903 10523
rect 25498 10520 25504 10532
rect 23891 10492 25504 10520
rect 23891 10489 23903 10492
rect 23845 10483 23903 10489
rect 25498 10480 25504 10492
rect 25556 10480 25562 10532
rect 28552 10520 28580 10560
rect 26353 10492 28580 10520
rect 20254 10452 20260 10464
rect 20215 10424 20260 10452
rect 20254 10412 20260 10424
rect 20312 10412 20318 10464
rect 20438 10412 20444 10464
rect 20496 10452 20502 10464
rect 26353 10452 26381 10492
rect 20496 10424 26381 10452
rect 20496 10412 20502 10424
rect 26418 10412 26424 10464
rect 26476 10452 26482 10464
rect 29917 10455 29975 10461
rect 29917 10452 29929 10455
rect 26476 10424 29929 10452
rect 26476 10412 26482 10424
rect 29917 10421 29929 10424
rect 29963 10421 29975 10455
rect 38010 10452 38016 10464
rect 37971 10424 38016 10452
rect 29917 10415 29975 10421
rect 38010 10412 38016 10424
rect 38068 10412 38074 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 15930 10248 15936 10260
rect 15891 10220 15936 10248
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 16485 10251 16543 10257
rect 16485 10217 16497 10251
rect 16531 10248 16543 10251
rect 16666 10248 16672 10260
rect 16531 10220 16672 10248
rect 16531 10217 16543 10220
rect 16485 10211 16543 10217
rect 15378 10112 15384 10124
rect 15339 10084 15384 10112
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 15473 10115 15531 10121
rect 15473 10081 15485 10115
rect 15519 10112 15531 10115
rect 16500 10112 16528 10211
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 18322 10248 18328 10260
rect 18283 10220 18328 10248
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 18506 10208 18512 10260
rect 18564 10248 18570 10260
rect 22462 10248 22468 10260
rect 18564 10220 22468 10248
rect 18564 10208 18570 10220
rect 22462 10208 22468 10220
rect 22520 10208 22526 10260
rect 27154 10208 27160 10260
rect 27212 10248 27218 10260
rect 27341 10251 27399 10257
rect 27341 10248 27353 10251
rect 27212 10220 27353 10248
rect 27212 10208 27218 10220
rect 27341 10217 27353 10220
rect 27387 10217 27399 10251
rect 27341 10211 27399 10217
rect 15519 10084 16528 10112
rect 17773 10115 17831 10121
rect 15519 10081 15531 10084
rect 15473 10075 15531 10081
rect 17773 10081 17785 10115
rect 17819 10112 17831 10115
rect 18230 10112 18236 10124
rect 17819 10084 18236 10112
rect 17819 10081 17831 10084
rect 17773 10075 17831 10081
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 20162 10112 20168 10124
rect 19904 10084 20168 10112
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 19794 10044 19800 10056
rect 19392 10016 19800 10044
rect 19392 10004 19398 10016
rect 19794 10004 19800 10016
rect 19852 10004 19858 10056
rect 19904 10053 19932 10084
rect 20162 10072 20168 10084
rect 20220 10072 20226 10124
rect 23198 10112 23204 10124
rect 23159 10084 23204 10112
rect 23198 10072 23204 10084
rect 23256 10072 23262 10124
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10013 19947 10047
rect 19889 10007 19947 10013
rect 20073 10047 20131 10053
rect 20073 10013 20085 10047
rect 20119 10044 20131 10047
rect 20533 10047 20591 10053
rect 20533 10044 20545 10047
rect 20119 10016 20545 10044
rect 20119 10013 20131 10016
rect 20073 10007 20131 10013
rect 20533 10013 20545 10016
rect 20579 10013 20591 10047
rect 26050 10044 26056 10056
rect 26011 10016 26056 10044
rect 20533 10007 20591 10013
rect 26050 10004 26056 10016
rect 26108 10044 26114 10056
rect 30466 10044 30472 10056
rect 26108 10016 30472 10044
rect 26108 10004 26114 10016
rect 30466 10004 30472 10016
rect 30524 10044 30530 10056
rect 31205 10047 31263 10053
rect 31205 10044 31217 10047
rect 30524 10016 31217 10044
rect 30524 10004 30530 10016
rect 31205 10013 31217 10016
rect 31251 10044 31263 10047
rect 33778 10044 33784 10056
rect 31251 10016 33784 10044
rect 31251 10013 31263 10016
rect 31205 10007 31263 10013
rect 33778 10004 33784 10016
rect 33836 10004 33842 10056
rect 14550 9936 14556 9988
rect 14608 9976 14614 9988
rect 15565 9979 15623 9985
rect 15565 9976 15577 9979
rect 14608 9948 15577 9976
rect 14608 9936 14614 9948
rect 15565 9945 15577 9948
rect 15611 9945 15623 9979
rect 15565 9939 15623 9945
rect 17865 9979 17923 9985
rect 17865 9945 17877 9979
rect 17911 9976 17923 9979
rect 18506 9976 18512 9988
rect 17911 9948 18512 9976
rect 17911 9945 17923 9948
rect 17865 9939 17923 9945
rect 18506 9936 18512 9948
rect 18564 9936 18570 9988
rect 18598 9936 18604 9988
rect 18656 9976 18662 9988
rect 22934 9979 22992 9985
rect 22934 9976 22946 9979
rect 18656 9948 22946 9976
rect 18656 9936 18662 9948
rect 22934 9945 22946 9948
rect 22980 9945 22992 9979
rect 22934 9939 22992 9945
rect 16666 9868 16672 9920
rect 16724 9908 16730 9920
rect 17957 9911 18015 9917
rect 17957 9908 17969 9911
rect 16724 9880 17969 9908
rect 16724 9868 16730 9880
rect 17957 9877 17969 9880
rect 18003 9877 18015 9911
rect 17957 9871 18015 9877
rect 20717 9911 20775 9917
rect 20717 9877 20729 9911
rect 20763 9908 20775 9911
rect 21358 9908 21364 9920
rect 20763 9880 21364 9908
rect 20763 9877 20775 9880
rect 20717 9871 20775 9877
rect 21358 9868 21364 9880
rect 21416 9868 21422 9920
rect 21818 9908 21824 9920
rect 21779 9880 21824 9908
rect 21818 9868 21824 9880
rect 21876 9868 21882 9920
rect 23566 9868 23572 9920
rect 23624 9908 23630 9920
rect 23842 9908 23848 9920
rect 23624 9880 23848 9908
rect 23624 9868 23630 9880
rect 23842 9868 23848 9880
rect 23900 9868 23906 9920
rect 31938 9868 31944 9920
rect 31996 9908 32002 9920
rect 32493 9911 32551 9917
rect 32493 9908 32505 9911
rect 31996 9880 32505 9908
rect 31996 9868 32002 9880
rect 32493 9877 32505 9880
rect 32539 9877 32551 9911
rect 32493 9871 32551 9877
rect 37369 9911 37427 9917
rect 37369 9877 37381 9911
rect 37415 9908 37427 9911
rect 37642 9908 37648 9920
rect 37415 9880 37648 9908
rect 37415 9877 37427 9880
rect 37369 9871 37427 9877
rect 37642 9868 37648 9880
rect 37700 9868 37706 9920
rect 37826 9908 37832 9920
rect 37787 9880 37832 9908
rect 37826 9868 37832 9880
rect 37884 9868 37890 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 11514 9704 11520 9716
rect 11475 9676 11520 9704
rect 11514 9664 11520 9676
rect 11572 9664 11578 9716
rect 18506 9704 18512 9716
rect 18467 9676 18512 9704
rect 18506 9664 18512 9676
rect 18564 9664 18570 9716
rect 20901 9707 20959 9713
rect 20901 9673 20913 9707
rect 20947 9673 20959 9707
rect 20901 9667 20959 9673
rect 9030 9596 9036 9648
rect 9088 9636 9094 9648
rect 10226 9636 10232 9648
rect 9088 9608 10232 9636
rect 9088 9596 9094 9608
rect 10226 9596 10232 9608
rect 10284 9636 10290 9648
rect 10781 9639 10839 9645
rect 10781 9636 10793 9639
rect 10284 9608 10793 9636
rect 10284 9596 10290 9608
rect 10781 9605 10793 9608
rect 10827 9605 10839 9639
rect 11974 9636 11980 9648
rect 11935 9608 11980 9636
rect 10781 9599 10839 9605
rect 11974 9596 11980 9608
rect 12032 9636 12038 9648
rect 14369 9639 14427 9645
rect 12032 9608 12434 9636
rect 12032 9596 12038 9608
rect 5810 9528 5816 9580
rect 5868 9568 5874 9580
rect 11885 9571 11943 9577
rect 11885 9568 11897 9571
rect 5868 9540 11897 9568
rect 5868 9528 5874 9540
rect 11885 9537 11897 9540
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 11974 9460 11980 9512
rect 12032 9500 12038 9512
rect 12069 9503 12127 9509
rect 12069 9500 12081 9503
rect 12032 9472 12081 9500
rect 12032 9460 12038 9472
rect 12069 9469 12081 9472
rect 12115 9469 12127 9503
rect 12406 9500 12434 9608
rect 14369 9605 14381 9639
rect 14415 9636 14427 9639
rect 15197 9639 15255 9645
rect 15197 9636 15209 9639
rect 14415 9608 15209 9636
rect 14415 9605 14427 9608
rect 14369 9599 14427 9605
rect 15197 9605 15209 9608
rect 15243 9636 15255 9639
rect 15286 9636 15292 9648
rect 15243 9608 15292 9636
rect 15243 9605 15255 9608
rect 15197 9599 15255 9605
rect 15286 9596 15292 9608
rect 15344 9596 15350 9648
rect 17770 9596 17776 9648
rect 17828 9636 17834 9648
rect 17828 9608 19104 9636
rect 17828 9596 17834 9608
rect 13446 9528 13452 9580
rect 13504 9568 13510 9580
rect 19076 9577 19104 9608
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 13504 9540 14289 9568
rect 13504 9528 13510 9540
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 19061 9571 19119 9577
rect 19061 9537 19073 9571
rect 19107 9537 19119 9571
rect 19061 9531 19119 9537
rect 19245 9571 19303 9577
rect 19245 9537 19257 9571
rect 19291 9568 19303 9571
rect 19334 9568 19340 9580
rect 19291 9540 19340 9568
rect 19291 9537 19303 9540
rect 19245 9531 19303 9537
rect 12802 9500 12808 9512
rect 12406 9472 12808 9500
rect 12069 9463 12127 9469
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 14553 9503 14611 9509
rect 14553 9469 14565 9503
rect 14599 9500 14611 9503
rect 15378 9500 15384 9512
rect 14599 9472 15384 9500
rect 14599 9469 14611 9472
rect 14553 9463 14611 9469
rect 15378 9460 15384 9472
rect 15436 9460 15442 9512
rect 16761 9503 16819 9509
rect 16761 9500 16773 9503
rect 16040 9472 16773 9500
rect 13354 9392 13360 9444
rect 13412 9432 13418 9444
rect 13909 9435 13967 9441
rect 13909 9432 13921 9435
rect 13412 9404 13921 9432
rect 13412 9392 13418 9404
rect 13909 9401 13921 9404
rect 13955 9401 13967 9435
rect 13909 9395 13967 9401
rect 14458 9324 14464 9376
rect 14516 9364 14522 9376
rect 16040 9373 16068 9472
rect 16761 9469 16773 9472
rect 16807 9469 16819 9503
rect 16868 9500 16896 9531
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 19429 9571 19487 9577
rect 19429 9537 19441 9571
rect 19475 9568 19487 9571
rect 20073 9571 20131 9577
rect 20073 9568 20085 9571
rect 19475 9540 20085 9568
rect 19475 9537 19487 9540
rect 19429 9531 19487 9537
rect 20073 9537 20085 9540
rect 20119 9537 20131 9571
rect 20714 9568 20720 9580
rect 20675 9540 20720 9568
rect 20073 9531 20131 9537
rect 20714 9528 20720 9540
rect 20772 9528 20778 9580
rect 17770 9500 17776 9512
rect 16868 9472 17776 9500
rect 16761 9463 16819 9469
rect 16776 9432 16804 9463
rect 17770 9460 17776 9472
rect 17828 9460 17834 9512
rect 20916 9500 20944 9667
rect 21358 9664 21364 9716
rect 21416 9704 21422 9716
rect 30558 9704 30564 9716
rect 21416 9676 30564 9704
rect 21416 9664 21422 9676
rect 30558 9664 30564 9676
rect 30616 9664 30622 9716
rect 23198 9636 23204 9648
rect 22204 9608 23204 9636
rect 22204 9577 22232 9608
rect 23198 9596 23204 9608
rect 23256 9596 23262 9648
rect 23382 9596 23388 9648
rect 23440 9636 23446 9648
rect 25142 9639 25200 9645
rect 25142 9636 25154 9639
rect 23440 9608 25154 9636
rect 23440 9596 23446 9608
rect 25142 9605 25154 9608
rect 25188 9605 25200 9639
rect 30386 9639 30444 9645
rect 30386 9636 30398 9639
rect 25142 9599 25200 9605
rect 25240 9608 30398 9636
rect 22189 9571 22247 9577
rect 22189 9537 22201 9571
rect 22235 9537 22247 9571
rect 22445 9571 22503 9577
rect 22445 9568 22457 9571
rect 22189 9531 22247 9537
rect 22296 9540 22457 9568
rect 20916 9472 21496 9500
rect 18690 9432 18696 9444
rect 16776 9404 18696 9432
rect 18690 9392 18696 9404
rect 18748 9392 18754 9444
rect 20257 9435 20315 9441
rect 20257 9401 20269 9435
rect 20303 9432 20315 9435
rect 21468 9432 21496 9472
rect 21542 9460 21548 9512
rect 21600 9500 21606 9512
rect 22296 9500 22324 9540
rect 22445 9537 22457 9540
rect 22491 9537 22503 9571
rect 25240 9568 25268 9608
rect 30386 9605 30398 9608
rect 30432 9605 30444 9639
rect 34158 9639 34216 9645
rect 34158 9636 34170 9639
rect 30386 9599 30444 9605
rect 30484 9608 34170 9636
rect 22445 9531 22503 9537
rect 23492 9540 25268 9568
rect 25409 9571 25467 9577
rect 21600 9472 22324 9500
rect 21600 9460 21606 9472
rect 22186 9432 22192 9444
rect 20303 9404 21220 9432
rect 21468 9404 22192 9432
rect 20303 9401 20315 9404
rect 20257 9395 20315 9401
rect 16025 9367 16083 9373
rect 16025 9364 16037 9367
rect 14516 9336 16037 9364
rect 14516 9324 14522 9336
rect 16025 9333 16037 9336
rect 16071 9333 16083 9367
rect 16025 9327 16083 9333
rect 17221 9367 17279 9373
rect 17221 9333 17233 9367
rect 17267 9364 17279 9367
rect 17494 9364 17500 9376
rect 17267 9336 17500 9364
rect 17267 9333 17279 9336
rect 17221 9327 17279 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 17770 9364 17776 9376
rect 17731 9336 17776 9364
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 21192 9364 21220 9404
rect 22186 9392 22192 9404
rect 22244 9392 22250 9444
rect 23492 9364 23520 9540
rect 25409 9537 25421 9571
rect 25455 9568 25467 9571
rect 25498 9568 25504 9580
rect 25455 9540 25504 9568
rect 25455 9537 25467 9540
rect 25409 9531 25467 9537
rect 25498 9528 25504 9540
rect 25556 9528 25562 9580
rect 28086 9571 28144 9577
rect 28086 9568 28098 9571
rect 25608 9540 28098 9568
rect 23566 9392 23572 9444
rect 23624 9432 23630 9444
rect 23624 9404 23669 9432
rect 23624 9392 23630 9404
rect 24026 9364 24032 9376
rect 21192 9336 23520 9364
rect 23987 9336 24032 9364
rect 24026 9324 24032 9336
rect 24084 9324 24090 9376
rect 24762 9324 24768 9376
rect 24820 9364 24826 9376
rect 25608 9364 25636 9540
rect 28086 9537 28098 9540
rect 28132 9537 28144 9571
rect 28350 9568 28356 9580
rect 28311 9540 28356 9568
rect 28086 9531 28144 9537
rect 28350 9528 28356 9540
rect 28408 9528 28414 9580
rect 30484 9568 30512 9608
rect 34158 9605 34170 9608
rect 34204 9605 34216 9639
rect 35526 9636 35532 9648
rect 34158 9599 34216 9605
rect 34900 9608 35532 9636
rect 28460 9540 30512 9568
rect 30653 9571 30711 9577
rect 26970 9364 26976 9376
rect 24820 9336 25636 9364
rect 26931 9336 26976 9364
rect 24820 9324 24826 9336
rect 26970 9324 26976 9336
rect 27028 9324 27034 9376
rect 27430 9324 27436 9376
rect 27488 9364 27494 9376
rect 28460 9364 28488 9540
rect 30653 9537 30665 9571
rect 30699 9568 30711 9571
rect 31938 9568 31944 9580
rect 30699 9540 31944 9568
rect 30699 9537 30711 9540
rect 30653 9531 30711 9537
rect 31938 9528 31944 9540
rect 31996 9528 32002 9580
rect 34900 9577 34928 9608
rect 35526 9596 35532 9608
rect 35584 9596 35590 9648
rect 34425 9571 34483 9577
rect 34425 9537 34437 9571
rect 34471 9568 34483 9571
rect 34885 9571 34943 9577
rect 34885 9568 34897 9571
rect 34471 9540 34897 9568
rect 34471 9537 34483 9540
rect 34425 9531 34483 9537
rect 34885 9537 34897 9540
rect 34931 9537 34943 9571
rect 35141 9571 35199 9577
rect 35141 9568 35153 9571
rect 34885 9531 34943 9537
rect 34992 9540 35153 9568
rect 34790 9460 34796 9512
rect 34848 9500 34854 9512
rect 34992 9500 35020 9540
rect 35141 9537 35153 9540
rect 35187 9537 35199 9571
rect 35141 9531 35199 9537
rect 34848 9472 35020 9500
rect 34848 9460 34854 9472
rect 29270 9364 29276 9376
rect 27488 9336 28488 9364
rect 29231 9336 29276 9364
rect 27488 9324 27494 9336
rect 29270 9324 29276 9336
rect 29328 9324 29334 9376
rect 29362 9324 29368 9376
rect 29420 9364 29426 9376
rect 33045 9367 33103 9373
rect 33045 9364 33057 9367
rect 29420 9336 33057 9364
rect 29420 9324 29426 9336
rect 33045 9333 33057 9336
rect 33091 9333 33103 9367
rect 33045 9327 33103 9333
rect 35618 9324 35624 9376
rect 35676 9364 35682 9376
rect 36265 9367 36323 9373
rect 36265 9364 36277 9367
rect 35676 9336 36277 9364
rect 35676 9324 35682 9336
rect 36265 9333 36277 9336
rect 36311 9333 36323 9367
rect 37734 9364 37740 9376
rect 37695 9336 37740 9364
rect 36265 9327 36323 9333
rect 37734 9324 37740 9336
rect 37792 9324 37798 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 14277 9163 14335 9169
rect 14277 9129 14289 9163
rect 14323 9160 14335 9163
rect 18598 9160 18604 9172
rect 14323 9132 18604 9160
rect 14323 9129 14335 9132
rect 14277 9123 14335 9129
rect 18598 9120 18604 9132
rect 18656 9120 18662 9172
rect 18690 9120 18696 9172
rect 18748 9160 18754 9172
rect 19981 9163 20039 9169
rect 18748 9132 18793 9160
rect 18748 9120 18754 9132
rect 19981 9129 19993 9163
rect 20027 9160 20039 9163
rect 20714 9160 20720 9172
rect 20027 9132 20720 9160
rect 20027 9129 20039 9132
rect 19981 9123 20039 9129
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 26418 9160 26424 9172
rect 21652 9132 26280 9160
rect 26379 9132 26424 9160
rect 10410 9092 10416 9104
rect 10060 9064 10416 9092
rect 10060 9033 10088 9064
rect 10410 9052 10416 9064
rect 10468 9092 10474 9104
rect 11974 9092 11980 9104
rect 10468 9064 11980 9092
rect 10468 9052 10474 9064
rect 11974 9052 11980 9064
rect 12032 9052 12038 9104
rect 14826 9092 14832 9104
rect 14787 9064 14832 9092
rect 14826 9052 14832 9064
rect 14884 9052 14890 9104
rect 17497 9095 17555 9101
rect 17497 9061 17509 9095
rect 17543 9092 17555 9095
rect 21542 9092 21548 9104
rect 17543 9064 21548 9092
rect 17543 9061 17555 9064
rect 17497 9055 17555 9061
rect 21542 9052 21548 9064
rect 21600 9052 21606 9104
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 8993 10103 9027
rect 10226 9024 10232 9036
rect 10187 8996 10232 9024
rect 10045 8987 10103 8993
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 12434 9024 12440 9036
rect 12406 8984 12440 9024
rect 12492 9024 12498 9036
rect 16945 9027 17003 9033
rect 16945 9024 16957 9027
rect 12492 8996 16957 9024
rect 12492 8984 12498 8996
rect 16945 8993 16957 8996
rect 16991 9024 17003 9027
rect 16991 8996 17724 9024
rect 16991 8993 17003 8996
rect 16945 8987 17003 8993
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8956 11667 8959
rect 12253 8959 12311 8965
rect 12253 8956 12265 8959
rect 11655 8928 12265 8956
rect 11655 8925 11667 8928
rect 11609 8919 11667 8925
rect 12253 8925 12265 8928
rect 12299 8956 12311 8959
rect 12406 8956 12434 8984
rect 12299 8928 12434 8956
rect 12299 8925 12311 8928
rect 12253 8919 12311 8925
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13964 8928 14105 8956
rect 13964 8916 13970 8928
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 17494 8956 17500 8968
rect 17455 8928 17500 8956
rect 14093 8919 14151 8925
rect 17494 8916 17500 8928
rect 17552 8916 17558 8968
rect 17696 8965 17724 8996
rect 18690 8984 18696 9036
rect 18748 9024 18754 9036
rect 19334 9024 19340 9036
rect 18748 8996 19340 9024
rect 18748 8984 18754 8996
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 19521 9027 19579 9033
rect 19521 8993 19533 9027
rect 19567 9024 19579 9027
rect 20530 9024 20536 9036
rect 19567 8996 20536 9024
rect 19567 8993 19579 8996
rect 19521 8987 19579 8993
rect 20530 8984 20536 8996
rect 20588 8984 20594 9036
rect 17681 8959 17739 8965
rect 17681 8925 17693 8959
rect 17727 8925 17739 8959
rect 17681 8919 17739 8925
rect 17862 8916 17868 8968
rect 17920 8956 17926 8968
rect 21652 8956 21680 9132
rect 26252 9092 26280 9132
rect 26418 9120 26424 9132
rect 26476 9120 26482 9172
rect 27338 9120 27344 9172
rect 27396 9160 27402 9172
rect 27433 9163 27491 9169
rect 27433 9160 27445 9163
rect 27396 9132 27445 9160
rect 27396 9120 27402 9132
rect 27433 9129 27445 9132
rect 27479 9129 27491 9163
rect 29178 9160 29184 9172
rect 27433 9123 27491 9129
rect 27908 9132 29184 9160
rect 27908 9092 27936 9132
rect 29178 9120 29184 9132
rect 29236 9120 29242 9172
rect 30561 9163 30619 9169
rect 30561 9129 30573 9163
rect 30607 9160 30619 9163
rect 30650 9160 30656 9172
rect 30607 9132 30656 9160
rect 30607 9129 30619 9132
rect 30561 9123 30619 9129
rect 30650 9120 30656 9132
rect 30708 9120 30714 9172
rect 33226 9160 33232 9172
rect 33187 9132 33232 9160
rect 33226 9120 33232 9132
rect 33284 9120 33290 9172
rect 34790 9120 34796 9172
rect 34848 9160 34854 9172
rect 34885 9163 34943 9169
rect 34885 9160 34897 9163
rect 34848 9132 34897 9160
rect 34848 9120 34854 9132
rect 34885 9129 34897 9132
rect 34931 9129 34943 9163
rect 34885 9123 34943 9129
rect 26252 9064 27936 9092
rect 33594 9052 33600 9104
rect 33652 9092 33658 9104
rect 34330 9092 34336 9104
rect 33652 9064 34336 9092
rect 33652 9052 33658 9064
rect 34330 9052 34336 9064
rect 34388 9092 34394 9104
rect 35621 9095 35679 9101
rect 35621 9092 35633 9095
rect 34388 9064 35633 9092
rect 34388 9052 34394 9064
rect 35621 9061 35633 9064
rect 35667 9061 35679 9095
rect 35621 9055 35679 9061
rect 22925 9027 22983 9033
rect 22925 8993 22937 9027
rect 22971 9024 22983 9027
rect 23198 9024 23204 9036
rect 22971 8996 23204 9024
rect 22971 8993 22983 8996
rect 22925 8987 22983 8993
rect 23198 8984 23204 8996
rect 23256 8984 23262 9036
rect 17920 8928 21680 8956
rect 25066 8959 25124 8965
rect 17920 8916 17926 8928
rect 25066 8925 25078 8959
rect 25112 8956 25124 8959
rect 28813 8959 28871 8965
rect 28813 8956 28825 8959
rect 25112 8928 25544 8956
rect 25112 8925 25124 8928
rect 25066 8919 25124 8925
rect 25516 8900 25544 8928
rect 28368 8928 28825 8956
rect 28368 8900 28396 8928
rect 28813 8925 28825 8928
rect 28859 8925 28871 8959
rect 28813 8919 28871 8925
rect 30558 8916 30564 8968
rect 30616 8956 30622 8968
rect 31674 8959 31732 8965
rect 31674 8956 31686 8959
rect 30616 8928 31686 8956
rect 30616 8916 30622 8928
rect 31674 8925 31686 8928
rect 31720 8925 31732 8959
rect 31938 8956 31944 8968
rect 31851 8928 31944 8956
rect 31674 8919 31732 8925
rect 31938 8916 31944 8928
rect 31996 8956 32002 8968
rect 32398 8956 32404 8968
rect 31996 8928 32404 8956
rect 31996 8916 32002 8928
rect 32398 8916 32404 8928
rect 32456 8916 32462 8968
rect 34698 8956 34704 8968
rect 34659 8928 34704 8956
rect 34698 8916 34704 8928
rect 34756 8916 34762 8968
rect 35526 8916 35532 8968
rect 35584 8956 35590 8968
rect 37001 8959 37059 8965
rect 37001 8956 37013 8959
rect 35584 8928 37013 8956
rect 35584 8916 35590 8928
rect 37001 8925 37013 8928
rect 37047 8925 37059 8959
rect 37001 8919 37059 8925
rect 9858 8848 9864 8900
rect 9916 8888 9922 8900
rect 10321 8891 10379 8897
rect 10321 8888 10333 8891
rect 9916 8860 10333 8888
rect 9916 8848 9922 8860
rect 10321 8857 10333 8860
rect 10367 8857 10379 8891
rect 10321 8851 10379 8857
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 13320 8860 15700 8888
rect 13320 8848 13326 8860
rect 10686 8820 10692 8832
rect 10647 8792 10692 8820
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 10962 8780 10968 8832
rect 11020 8820 11026 8832
rect 11701 8823 11759 8829
rect 11701 8820 11713 8823
rect 11020 8792 11713 8820
rect 11020 8780 11026 8792
rect 11701 8789 11713 8792
rect 11747 8820 11759 8823
rect 15562 8820 15568 8832
rect 11747 8792 15568 8820
rect 11747 8789 11759 8792
rect 11701 8783 11759 8789
rect 15562 8780 15568 8792
rect 15620 8780 15626 8832
rect 15672 8820 15700 8860
rect 17770 8848 17776 8900
rect 17828 8888 17834 8900
rect 17828 8860 21680 8888
rect 17828 8848 17834 8860
rect 19613 8823 19671 8829
rect 19613 8820 19625 8823
rect 15672 8792 19625 8820
rect 19613 8789 19625 8792
rect 19659 8820 19671 8823
rect 20993 8823 21051 8829
rect 20993 8820 21005 8823
rect 19659 8792 21005 8820
rect 19659 8789 19671 8792
rect 19613 8783 19671 8789
rect 20993 8789 21005 8792
rect 21039 8789 21051 8823
rect 20993 8783 21051 8789
rect 21082 8780 21088 8832
rect 21140 8820 21146 8832
rect 21545 8823 21603 8829
rect 21545 8820 21557 8823
rect 21140 8792 21557 8820
rect 21140 8780 21146 8792
rect 21545 8789 21557 8792
rect 21591 8789 21603 8823
rect 21652 8820 21680 8860
rect 21726 8848 21732 8900
rect 21784 8888 21790 8900
rect 22658 8891 22716 8897
rect 22658 8888 22670 8891
rect 21784 8860 22670 8888
rect 21784 8848 21790 8860
rect 22658 8857 22670 8860
rect 22704 8857 22716 8891
rect 22658 8851 22716 8857
rect 22830 8848 22836 8900
rect 22888 8888 22894 8900
rect 22888 8860 24817 8888
rect 22888 8848 22894 8860
rect 23566 8820 23572 8832
rect 21652 8792 23572 8820
rect 21545 8783 21603 8789
rect 23566 8780 23572 8792
rect 23624 8780 23630 8832
rect 24789 8820 24817 8860
rect 24854 8848 24860 8900
rect 24912 8888 24918 8900
rect 25286 8891 25344 8897
rect 25286 8888 25298 8891
rect 24912 8860 25298 8888
rect 24912 8848 24918 8860
rect 25286 8857 25298 8860
rect 25332 8857 25344 8891
rect 25286 8851 25344 8857
rect 25498 8848 25504 8900
rect 25556 8848 25562 8900
rect 26326 8848 26332 8900
rect 26384 8888 26390 8900
rect 26384 8860 27568 8888
rect 26384 8848 26390 8860
rect 26970 8820 26976 8832
rect 24789 8792 26976 8820
rect 26970 8780 26976 8792
rect 27028 8780 27034 8832
rect 27540 8820 27568 8860
rect 28350 8848 28356 8900
rect 28408 8848 28414 8900
rect 28546 8891 28604 8897
rect 28546 8888 28558 8891
rect 28460 8860 28558 8888
rect 28460 8820 28488 8860
rect 28546 8857 28558 8860
rect 28592 8857 28604 8891
rect 28546 8851 28604 8857
rect 34146 8848 34152 8900
rect 34204 8888 34210 8900
rect 36734 8891 36792 8897
rect 36734 8888 36746 8891
rect 34204 8860 36746 8888
rect 34204 8848 34210 8860
rect 36734 8857 36746 8860
rect 36780 8857 36792 8891
rect 36734 8851 36792 8857
rect 27540 8792 28488 8820
rect 33873 8823 33931 8829
rect 33873 8789 33885 8823
rect 33919 8820 33931 8823
rect 34054 8820 34060 8832
rect 33919 8792 34060 8820
rect 33919 8789 33931 8792
rect 33873 8783 33931 8789
rect 34054 8780 34060 8792
rect 34112 8780 34118 8832
rect 36998 8780 37004 8832
rect 37056 8820 37062 8832
rect 37461 8823 37519 8829
rect 37461 8820 37473 8823
rect 37056 8792 37473 8820
rect 37056 8780 37062 8792
rect 37461 8789 37473 8792
rect 37507 8789 37519 8823
rect 37461 8783 37519 8789
rect 37918 8780 37924 8832
rect 37976 8820 37982 8832
rect 38013 8823 38071 8829
rect 38013 8820 38025 8823
rect 37976 8792 38025 8820
rect 37976 8780 37982 8792
rect 38013 8789 38025 8792
rect 38059 8789 38071 8823
rect 38013 8783 38071 8789
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 10870 8616 10876 8628
rect 10831 8588 10876 8616
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 11977 8619 12035 8625
rect 11977 8585 11989 8619
rect 12023 8616 12035 8619
rect 12618 8616 12624 8628
rect 12023 8588 12624 8616
rect 12023 8585 12035 8588
rect 11977 8579 12035 8585
rect 12618 8576 12624 8588
rect 12676 8616 12682 8628
rect 13722 8616 13728 8628
rect 12676 8588 13728 8616
rect 12676 8576 12682 8588
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 13906 8616 13912 8628
rect 13867 8588 13912 8616
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 14369 8619 14427 8625
rect 14369 8585 14381 8619
rect 14415 8616 14427 8619
rect 14826 8616 14832 8628
rect 14415 8588 14832 8616
rect 14415 8585 14427 8588
rect 14369 8579 14427 8585
rect 14826 8576 14832 8588
rect 14884 8576 14890 8628
rect 15378 8576 15384 8628
rect 15436 8576 15442 8628
rect 15930 8616 15936 8628
rect 15843 8588 15936 8616
rect 15930 8576 15936 8588
rect 15988 8616 15994 8628
rect 16390 8616 16396 8628
rect 15988 8588 16396 8616
rect 15988 8576 15994 8588
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 20070 8576 20076 8628
rect 20128 8616 20134 8628
rect 29270 8616 29276 8628
rect 20128 8588 21036 8616
rect 20128 8576 20134 8588
rect 8662 8508 8668 8560
rect 8720 8548 8726 8560
rect 12069 8551 12127 8557
rect 12069 8548 12081 8551
rect 8720 8520 12081 8548
rect 8720 8508 8726 8520
rect 12069 8517 12081 8520
rect 12115 8517 12127 8551
rect 15396 8548 15424 8576
rect 16482 8548 16488 8560
rect 12069 8511 12127 8517
rect 14568 8520 16488 8548
rect 10686 8480 10692 8492
rect 10647 8452 10692 8480
rect 10686 8440 10692 8452
rect 10744 8440 10750 8492
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 12452 8452 13185 8480
rect 11885 8415 11943 8421
rect 11885 8381 11897 8415
rect 11931 8412 11943 8415
rect 11974 8412 11980 8424
rect 11931 8384 11980 8412
rect 11931 8381 11943 8384
rect 11885 8375 11943 8381
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 12452 8353 12480 8452
rect 13173 8449 13185 8452
rect 13219 8449 13231 8483
rect 14274 8480 14280 8492
rect 14235 8452 14280 8480
rect 13173 8443 13231 8449
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 14568 8421 14596 8520
rect 16482 8508 16488 8520
rect 16540 8508 16546 8560
rect 17954 8508 17960 8560
rect 18012 8508 18018 8560
rect 20438 8548 20444 8560
rect 19306 8520 20208 8548
rect 20399 8520 20444 8548
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8480 15255 8483
rect 15286 8480 15292 8492
rect 15243 8452 15292 8480
rect 15243 8449 15255 8452
rect 15197 8443 15255 8449
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8480 15439 8483
rect 15930 8480 15936 8492
rect 15427 8452 15936 8480
rect 15427 8449 15439 8452
rect 15381 8443 15439 8449
rect 15930 8440 15936 8452
rect 15988 8440 15994 8492
rect 18049 8483 18107 8489
rect 18049 8480 18061 8483
rect 17696 8452 18061 8480
rect 17696 8424 17724 8452
rect 18049 8449 18061 8452
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8480 18659 8483
rect 19306 8480 19334 8520
rect 18647 8452 19334 8480
rect 20180 8480 20208 8520
rect 20438 8508 20444 8520
rect 20496 8508 20502 8560
rect 21008 8557 21036 8588
rect 22112 8588 29276 8616
rect 20993 8551 21051 8557
rect 20993 8517 21005 8551
rect 21039 8548 21051 8551
rect 22002 8548 22008 8560
rect 21039 8520 22008 8548
rect 21039 8517 21051 8520
rect 20993 8511 21051 8517
rect 22002 8508 22008 8520
rect 22060 8508 22066 8560
rect 22112 8480 22140 8588
rect 29270 8576 29276 8588
rect 29328 8576 29334 8628
rect 34146 8616 34152 8628
rect 34107 8588 34152 8616
rect 34146 8576 34152 8588
rect 34204 8576 34210 8628
rect 35434 8576 35440 8628
rect 35492 8616 35498 8628
rect 36265 8619 36323 8625
rect 36265 8616 36277 8619
rect 35492 8588 36277 8616
rect 35492 8576 35498 8588
rect 36265 8585 36277 8588
rect 36311 8585 36323 8619
rect 36265 8579 36323 8585
rect 34606 8548 34612 8560
rect 22296 8520 34612 8548
rect 22296 8480 22324 8520
rect 34606 8508 34612 8520
rect 34664 8508 34670 8560
rect 35802 8548 35808 8560
rect 35763 8520 35808 8548
rect 35802 8508 35808 8520
rect 35860 8508 35866 8560
rect 20180 8452 22140 8480
rect 22204 8452 22324 8480
rect 18647 8449 18659 8452
rect 18601 8443 18659 8449
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8381 14611 8415
rect 14553 8375 14611 8381
rect 17678 8372 17684 8424
rect 17736 8372 17742 8424
rect 19797 8415 19855 8421
rect 19797 8381 19809 8415
rect 19843 8412 19855 8415
rect 19978 8412 19984 8424
rect 19843 8384 19984 8412
rect 19843 8381 19855 8384
rect 19797 8375 19855 8381
rect 19978 8372 19984 8384
rect 20036 8372 20042 8424
rect 20070 8372 20076 8424
rect 20128 8412 20134 8424
rect 20165 8415 20223 8421
rect 20165 8412 20177 8415
rect 20128 8384 20177 8412
rect 20128 8372 20134 8384
rect 20165 8381 20177 8384
rect 20211 8381 20223 8415
rect 20165 8375 20223 8381
rect 20257 8415 20315 8421
rect 20257 8381 20269 8415
rect 20303 8412 20315 8415
rect 20438 8412 20444 8424
rect 20303 8384 20444 8412
rect 20303 8381 20315 8384
rect 20257 8375 20315 8381
rect 20438 8372 20444 8384
rect 20496 8372 20502 8424
rect 21082 8372 21088 8424
rect 21140 8412 21146 8424
rect 21266 8412 21272 8424
rect 21140 8384 21272 8412
rect 21140 8372 21146 8384
rect 21266 8372 21272 8384
rect 21324 8412 21330 8424
rect 22204 8412 22232 8452
rect 22370 8440 22376 8492
rect 22428 8480 22434 8492
rect 22934 8483 22992 8489
rect 22934 8480 22946 8483
rect 22428 8452 22946 8480
rect 22428 8440 22434 8452
rect 22934 8449 22946 8452
rect 22980 8449 22992 8483
rect 23198 8480 23204 8492
rect 23159 8452 23204 8480
rect 22934 8443 22992 8449
rect 23198 8440 23204 8452
rect 23256 8440 23262 8492
rect 26234 8440 26240 8492
rect 26292 8480 26298 8492
rect 28086 8483 28144 8489
rect 28086 8480 28098 8483
rect 26292 8452 28098 8480
rect 26292 8440 26298 8452
rect 28086 8449 28098 8452
rect 28132 8449 28144 8483
rect 28350 8480 28356 8492
rect 28311 8452 28356 8480
rect 28086 8443 28144 8449
rect 28350 8440 28356 8452
rect 28408 8440 28414 8492
rect 33965 8483 34023 8489
rect 33965 8449 33977 8483
rect 34011 8480 34023 8483
rect 34422 8480 34428 8492
rect 34011 8452 34428 8480
rect 34011 8449 34023 8452
rect 33965 8443 34023 8449
rect 34422 8440 34428 8452
rect 34480 8440 34486 8492
rect 21324 8384 21864 8412
rect 21324 8372 21330 8384
rect 12437 8347 12495 8353
rect 12437 8313 12449 8347
rect 12483 8313 12495 8347
rect 12437 8307 12495 8313
rect 13357 8347 13415 8353
rect 13357 8313 13369 8347
rect 13403 8344 13415 8347
rect 21726 8344 21732 8356
rect 13403 8316 21732 8344
rect 13403 8313 13415 8316
rect 13357 8307 13415 8313
rect 21726 8304 21732 8316
rect 21784 8304 21790 8356
rect 21836 8353 21864 8384
rect 22066 8384 22232 8412
rect 21821 8347 21879 8353
rect 21821 8313 21833 8347
rect 21867 8313 21879 8347
rect 22066 8344 22094 8384
rect 21821 8307 21879 8313
rect 21928 8316 22094 8344
rect 15289 8279 15347 8285
rect 15289 8245 15301 8279
rect 15335 8276 15347 8279
rect 15378 8276 15384 8288
rect 15335 8248 15384 8276
rect 15335 8245 15347 8248
rect 15289 8239 15347 8245
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 20438 8236 20444 8288
rect 20496 8276 20502 8288
rect 21928 8276 21956 8316
rect 26142 8304 26148 8356
rect 26200 8344 26206 8356
rect 26973 8347 27031 8353
rect 26973 8344 26985 8347
rect 26200 8316 26985 8344
rect 26200 8304 26206 8316
rect 26973 8313 26985 8316
rect 27019 8313 27031 8347
rect 30650 8344 30656 8356
rect 26973 8307 27031 8313
rect 28368 8316 30656 8344
rect 20496 8248 21956 8276
rect 20496 8236 20502 8248
rect 22002 8236 22008 8288
rect 22060 8276 22066 8288
rect 26160 8276 26188 8304
rect 22060 8248 26188 8276
rect 22060 8236 22066 8248
rect 27430 8236 27436 8288
rect 27488 8276 27494 8288
rect 28368 8276 28396 8316
rect 30650 8304 30656 8316
rect 30708 8304 30714 8356
rect 37366 8344 37372 8356
rect 37327 8316 37372 8344
rect 37366 8304 37372 8316
rect 37424 8304 37430 8356
rect 37921 8347 37979 8353
rect 37921 8313 37933 8347
rect 37967 8344 37979 8347
rect 38102 8344 38108 8356
rect 37967 8316 38108 8344
rect 37967 8313 37979 8316
rect 37921 8307 37979 8313
rect 38102 8304 38108 8316
rect 38160 8304 38166 8356
rect 32214 8276 32220 8288
rect 27488 8248 28396 8276
rect 32175 8248 32220 8276
rect 27488 8236 27494 8248
rect 32214 8236 32220 8248
rect 32272 8236 32278 8288
rect 33321 8279 33379 8285
rect 33321 8245 33333 8279
rect 33367 8276 33379 8279
rect 34609 8279 34667 8285
rect 34609 8276 34621 8279
rect 33367 8248 34621 8276
rect 33367 8245 33379 8248
rect 33321 8239 33379 8245
rect 34609 8245 34621 8248
rect 34655 8276 34667 8279
rect 35161 8279 35219 8285
rect 35161 8276 35173 8279
rect 34655 8248 35173 8276
rect 34655 8245 34667 8248
rect 34609 8239 34667 8245
rect 35161 8245 35173 8248
rect 35207 8276 35219 8279
rect 35342 8276 35348 8288
rect 35207 8248 35348 8276
rect 35207 8245 35219 8248
rect 35161 8239 35219 8245
rect 35342 8236 35348 8248
rect 35400 8236 35406 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 10318 8032 10324 8084
rect 10376 8072 10382 8084
rect 11057 8075 11115 8081
rect 11057 8072 11069 8075
rect 10376 8044 11069 8072
rect 10376 8032 10382 8044
rect 11057 8041 11069 8044
rect 11103 8041 11115 8075
rect 12618 8072 12624 8084
rect 12579 8044 12624 8072
rect 11057 8035 11115 8041
rect 11072 8004 11100 8035
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 18049 8075 18107 8081
rect 18049 8041 18061 8075
rect 18095 8072 18107 8075
rect 24854 8072 24860 8084
rect 18095 8044 24860 8072
rect 18095 8041 18107 8044
rect 18049 8035 18107 8041
rect 24854 8032 24860 8044
rect 24912 8032 24918 8084
rect 30466 8072 30472 8084
rect 30427 8044 30472 8072
rect 30466 8032 30472 8044
rect 30524 8032 30530 8084
rect 30834 8032 30840 8084
rect 30892 8072 30898 8084
rect 33962 8072 33968 8084
rect 30892 8044 33968 8072
rect 30892 8032 30898 8044
rect 33962 8032 33968 8044
rect 34020 8032 34026 8084
rect 34698 8072 34704 8084
rect 34659 8044 34704 8072
rect 34698 8032 34704 8044
rect 34756 8032 34762 8084
rect 37090 8032 37096 8084
rect 37148 8072 37154 8084
rect 38105 8075 38163 8081
rect 38105 8072 38117 8075
rect 37148 8044 38117 8072
rect 37148 8032 37154 8044
rect 38105 8041 38117 8044
rect 38151 8041 38163 8075
rect 38105 8035 38163 8041
rect 15102 8004 15108 8016
rect 11072 7976 15108 8004
rect 15102 7964 15108 7976
rect 15160 7964 15166 8016
rect 18693 8007 18751 8013
rect 18693 7973 18705 8007
rect 18739 8004 18751 8007
rect 35618 8004 35624 8016
rect 18739 7976 22094 8004
rect 18739 7973 18751 7976
rect 18693 7967 18751 7973
rect 11146 7896 11152 7948
rect 11204 7936 11210 7948
rect 16577 7939 16635 7945
rect 16577 7936 16589 7939
rect 11204 7908 16589 7936
rect 11204 7896 11210 7908
rect 15194 7868 15200 7880
rect 15155 7840 15200 7868
rect 15194 7828 15200 7840
rect 15252 7828 15258 7880
rect 15378 7868 15384 7880
rect 15339 7840 15384 7868
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 15948 7877 15976 7908
rect 16577 7905 16589 7908
rect 16623 7936 16635 7939
rect 17954 7936 17960 7948
rect 16623 7908 17960 7936
rect 16623 7905 16635 7908
rect 16577 7899 16635 7905
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 19334 7896 19340 7948
rect 19392 7936 19398 7948
rect 19889 7939 19947 7945
rect 19889 7936 19901 7939
rect 19392 7908 19901 7936
rect 19392 7896 19398 7908
rect 19889 7905 19901 7908
rect 19935 7936 19947 7939
rect 20438 7936 20444 7948
rect 19935 7908 20444 7936
rect 19935 7905 19947 7908
rect 19889 7899 19947 7905
rect 20438 7896 20444 7908
rect 20496 7896 20502 7948
rect 15933 7871 15991 7877
rect 15933 7837 15945 7871
rect 15979 7837 15991 7871
rect 15933 7831 15991 7837
rect 17402 7828 17408 7880
rect 17460 7868 17466 7880
rect 17865 7871 17923 7877
rect 17865 7868 17877 7871
rect 17460 7840 17877 7868
rect 17460 7828 17466 7840
rect 17865 7837 17877 7840
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 18509 7871 18567 7877
rect 18509 7837 18521 7871
rect 18555 7868 18567 7871
rect 18690 7868 18696 7880
rect 18555 7840 18696 7868
rect 18555 7837 18567 7840
rect 18509 7831 18567 7837
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 19242 7868 19248 7880
rect 19203 7840 19248 7868
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 22066 7868 22094 7976
rect 35176 7976 35624 8004
rect 32398 7936 32404 7948
rect 32359 7908 32404 7936
rect 32398 7896 32404 7908
rect 32456 7896 32462 7948
rect 35176 7945 35204 7976
rect 35618 7964 35624 7976
rect 35676 7964 35682 8016
rect 35161 7939 35219 7945
rect 35161 7905 35173 7939
rect 35207 7905 35219 7939
rect 35342 7936 35348 7948
rect 35303 7908 35348 7936
rect 35161 7899 35219 7905
rect 35342 7896 35348 7908
rect 35400 7896 35406 7948
rect 23109 7871 23167 7877
rect 22066 7840 22968 7868
rect 12066 7760 12072 7812
rect 12124 7800 12130 7812
rect 19334 7800 19340 7812
rect 12124 7772 19340 7800
rect 12124 7760 12130 7772
rect 19334 7760 19340 7772
rect 19392 7760 19398 7812
rect 19444 7772 21864 7800
rect 16025 7735 16083 7741
rect 16025 7701 16037 7735
rect 16071 7732 16083 7735
rect 17034 7732 17040 7744
rect 16071 7704 17040 7732
rect 16071 7701 16083 7704
rect 16025 7695 16083 7701
rect 17034 7692 17040 7704
rect 17092 7692 17098 7744
rect 19444 7741 19472 7772
rect 19429 7735 19487 7741
rect 19429 7701 19441 7735
rect 19475 7701 19487 7735
rect 19429 7695 19487 7701
rect 20806 7692 20812 7744
rect 20864 7732 20870 7744
rect 21729 7735 21787 7741
rect 21729 7732 21741 7735
rect 20864 7704 21741 7732
rect 20864 7692 20870 7704
rect 21729 7701 21741 7704
rect 21775 7701 21787 7735
rect 21836 7732 21864 7772
rect 22278 7760 22284 7812
rect 22336 7800 22342 7812
rect 22842 7803 22900 7809
rect 22842 7800 22854 7803
rect 22336 7772 22854 7800
rect 22336 7760 22342 7772
rect 22842 7769 22854 7772
rect 22888 7769 22900 7803
rect 22940 7800 22968 7840
rect 23109 7837 23121 7871
rect 23155 7868 23167 7871
rect 23474 7868 23480 7880
rect 23155 7840 23480 7868
rect 23155 7837 23167 7840
rect 23109 7831 23167 7837
rect 23474 7828 23480 7840
rect 23532 7828 23538 7880
rect 27614 7868 27620 7880
rect 27575 7840 27620 7868
rect 27614 7828 27620 7840
rect 27672 7828 27678 7880
rect 31941 7871 31999 7877
rect 31941 7837 31953 7871
rect 31987 7868 31999 7871
rect 32214 7868 32220 7880
rect 31987 7840 32220 7868
rect 31987 7837 31999 7840
rect 31941 7831 31999 7837
rect 32214 7828 32220 7840
rect 32272 7868 32278 7880
rect 32272 7840 34100 7868
rect 32272 7828 32278 7840
rect 27350 7803 27408 7809
rect 27350 7800 27362 7803
rect 22940 7772 27362 7800
rect 22842 7763 22900 7769
rect 27350 7769 27362 7772
rect 27396 7769 27408 7803
rect 27350 7763 27408 7769
rect 29086 7760 29092 7812
rect 29144 7800 29150 7812
rect 32646 7803 32704 7809
rect 32646 7800 32658 7803
rect 29144 7772 32658 7800
rect 29144 7760 29150 7772
rect 32646 7769 32658 7772
rect 32692 7769 32704 7803
rect 34072 7800 34100 7840
rect 34790 7828 34796 7880
rect 34848 7868 34854 7880
rect 36081 7871 36139 7877
rect 36081 7868 36093 7871
rect 34848 7840 36093 7868
rect 34848 7828 34854 7840
rect 36081 7837 36093 7840
rect 36127 7837 36139 7871
rect 36081 7831 36139 7837
rect 36170 7828 36176 7880
rect 36228 7868 36234 7880
rect 36725 7871 36783 7877
rect 36725 7868 36737 7871
rect 36228 7840 36737 7868
rect 36228 7828 36234 7840
rect 36725 7837 36737 7840
rect 36771 7837 36783 7871
rect 38194 7868 38200 7880
rect 36725 7831 36783 7837
rect 36832 7840 38200 7868
rect 36832 7800 36860 7840
rect 38194 7828 38200 7840
rect 38252 7828 38258 7880
rect 36981 7803 37039 7809
rect 36981 7800 36993 7803
rect 34072 7772 36860 7800
rect 36924 7772 36993 7800
rect 32646 7763 32704 7769
rect 23750 7732 23756 7744
rect 21836 7704 23756 7732
rect 21729 7695 21787 7701
rect 23750 7692 23756 7704
rect 23808 7692 23814 7744
rect 26234 7732 26240 7744
rect 26195 7704 26240 7732
rect 26234 7692 26240 7704
rect 26292 7692 26298 7744
rect 33134 7692 33140 7744
rect 33192 7732 33198 7744
rect 33781 7735 33839 7741
rect 33781 7732 33793 7735
rect 33192 7704 33793 7732
rect 33192 7692 33198 7704
rect 33781 7701 33793 7704
rect 33827 7701 33839 7735
rect 33781 7695 33839 7701
rect 35069 7735 35127 7741
rect 35069 7701 35081 7735
rect 35115 7732 35127 7735
rect 35802 7732 35808 7744
rect 35115 7704 35808 7732
rect 35115 7701 35127 7704
rect 35069 7695 35127 7701
rect 35802 7692 35808 7704
rect 35860 7692 35866 7744
rect 36265 7735 36323 7741
rect 36265 7701 36277 7735
rect 36311 7732 36323 7735
rect 36924 7732 36952 7772
rect 36981 7769 36993 7772
rect 37027 7769 37039 7803
rect 36981 7763 37039 7769
rect 36311 7704 36952 7732
rect 36311 7701 36323 7704
rect 36265 7695 36323 7701
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 10318 7488 10324 7540
rect 10376 7528 10382 7540
rect 10505 7531 10563 7537
rect 10505 7528 10517 7531
rect 10376 7500 10517 7528
rect 10376 7488 10382 7500
rect 10505 7497 10517 7500
rect 10551 7497 10563 7531
rect 12066 7528 12072 7540
rect 12027 7500 12072 7528
rect 10505 7491 10563 7497
rect 12066 7488 12072 7500
rect 12124 7488 12130 7540
rect 15194 7488 15200 7540
rect 15252 7528 15258 7540
rect 15565 7531 15623 7537
rect 15565 7528 15577 7531
rect 15252 7500 15577 7528
rect 15252 7488 15258 7500
rect 15565 7497 15577 7500
rect 15611 7497 15623 7531
rect 15565 7491 15623 7497
rect 15930 7488 15936 7540
rect 15988 7528 15994 7540
rect 16025 7531 16083 7537
rect 16025 7528 16037 7531
rect 15988 7500 16037 7528
rect 15988 7488 15994 7500
rect 16025 7497 16037 7500
rect 16071 7497 16083 7531
rect 16942 7528 16948 7540
rect 16903 7500 16948 7528
rect 16025 7491 16083 7497
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17402 7528 17408 7540
rect 17363 7500 17408 7528
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 18690 7528 18696 7540
rect 18651 7500 18696 7528
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 19613 7531 19671 7537
rect 19613 7497 19625 7531
rect 19659 7497 19671 7531
rect 19613 7491 19671 7497
rect 20165 7531 20223 7537
rect 20165 7497 20177 7531
rect 20211 7528 20223 7531
rect 20714 7528 20720 7540
rect 20211 7500 20720 7528
rect 20211 7497 20223 7500
rect 20165 7491 20223 7497
rect 7006 7420 7012 7472
rect 7064 7460 7070 7472
rect 10597 7463 10655 7469
rect 10597 7460 10609 7463
rect 7064 7432 10609 7460
rect 7064 7420 7070 7432
rect 10597 7429 10609 7432
rect 10643 7429 10655 7463
rect 15286 7460 15292 7472
rect 15199 7432 15292 7460
rect 10597 7423 10655 7429
rect 9585 7395 9643 7401
rect 9585 7361 9597 7395
rect 9631 7392 9643 7395
rect 9950 7392 9956 7404
rect 9631 7364 9956 7392
rect 9631 7361 9643 7364
rect 9585 7355 9643 7361
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7392 11943 7395
rect 12158 7392 12164 7404
rect 11931 7364 12164 7392
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 12158 7352 12164 7364
rect 12216 7352 12222 7404
rect 13538 7392 13544 7404
rect 13499 7364 13544 7392
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 13722 7392 13728 7404
rect 13683 7364 13728 7392
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 15212 7401 15240 7432
rect 15286 7420 15292 7432
rect 15344 7460 15350 7472
rect 19628 7460 19656 7491
rect 20714 7488 20720 7500
rect 20772 7528 20778 7540
rect 26234 7528 26240 7540
rect 20772 7500 26240 7528
rect 20772 7488 20778 7500
rect 26234 7488 26240 7500
rect 26292 7488 26298 7540
rect 29086 7528 29092 7540
rect 29047 7500 29092 7528
rect 29086 7488 29092 7500
rect 29144 7488 29150 7540
rect 29549 7531 29607 7537
rect 29549 7497 29561 7531
rect 29595 7497 29607 7531
rect 34790 7528 34796 7540
rect 34751 7500 34796 7528
rect 29549 7491 29607 7497
rect 24274 7463 24332 7469
rect 24274 7460 24286 7463
rect 15344 7432 18644 7460
rect 19628 7432 24286 7460
rect 15344 7420 15350 7432
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7361 15255 7395
rect 15197 7355 15255 7361
rect 15381 7395 15439 7401
rect 15381 7361 15393 7395
rect 15427 7361 15439 7395
rect 15381 7355 15439 7361
rect 10410 7324 10416 7336
rect 10371 7296 10416 7324
rect 10410 7284 10416 7296
rect 10468 7284 10474 7336
rect 12618 7284 12624 7336
rect 12676 7324 12682 7336
rect 14185 7327 14243 7333
rect 14185 7324 14197 7327
rect 12676 7296 14197 7324
rect 12676 7284 12682 7296
rect 14185 7293 14197 7296
rect 14231 7324 14243 7327
rect 14458 7324 14464 7336
rect 14231 7296 14464 7324
rect 14231 7293 14243 7296
rect 14185 7287 14243 7293
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 15396 7324 15424 7355
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 15528 7364 17049 7392
rect 15528 7352 15534 7364
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 18325 7395 18383 7401
rect 18325 7361 18337 7395
rect 18371 7392 18383 7395
rect 18506 7392 18512 7404
rect 18371 7364 18512 7392
rect 18371 7361 18383 7364
rect 18325 7355 18383 7361
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 15930 7324 15936 7336
rect 15396 7296 15936 7324
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 16482 7284 16488 7336
rect 16540 7324 16546 7336
rect 16761 7327 16819 7333
rect 16761 7324 16773 7327
rect 16540 7296 16773 7324
rect 16540 7284 16546 7296
rect 16761 7293 16773 7296
rect 16807 7293 16819 7327
rect 18138 7324 18144 7336
rect 18099 7296 18144 7324
rect 16761 7287 16819 7293
rect 18138 7284 18144 7296
rect 18196 7284 18202 7336
rect 18233 7327 18291 7333
rect 18233 7293 18245 7327
rect 18279 7293 18291 7327
rect 18616 7324 18644 7432
rect 24274 7429 24286 7432
rect 24320 7429 24332 7463
rect 29564 7460 29592 7491
rect 34790 7488 34796 7500
rect 34848 7488 34854 7540
rect 35345 7531 35403 7537
rect 35345 7497 35357 7531
rect 35391 7528 35403 7531
rect 37090 7528 37096 7540
rect 35391 7500 37096 7528
rect 35391 7497 35403 7500
rect 35345 7491 35403 7497
rect 24274 7423 24332 7429
rect 24412 7432 29592 7460
rect 19426 7392 19432 7404
rect 19387 7364 19432 7392
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 24412 7392 24440 7432
rect 30374 7420 30380 7472
rect 30432 7460 30438 7472
rect 30662 7463 30720 7469
rect 30662 7460 30674 7463
rect 30432 7432 30674 7460
rect 30432 7420 30438 7432
rect 30662 7429 30674 7432
rect 30708 7429 30720 7463
rect 30662 7423 30720 7429
rect 34333 7463 34391 7469
rect 34333 7429 34345 7463
rect 34379 7460 34391 7463
rect 35360 7460 35388 7491
rect 37090 7488 37096 7500
rect 37148 7488 37154 7540
rect 34379 7432 35388 7460
rect 36449 7463 36507 7469
rect 34379 7429 34391 7432
rect 34333 7423 34391 7429
rect 36449 7429 36461 7463
rect 36495 7460 36507 7463
rect 37274 7460 37280 7472
rect 36495 7432 37280 7460
rect 36495 7429 36507 7432
rect 36449 7423 36507 7429
rect 37274 7420 37280 7432
rect 37332 7420 37338 7472
rect 22066 7364 24440 7392
rect 28905 7395 28963 7401
rect 22066 7324 22094 7364
rect 28905 7361 28917 7395
rect 28951 7392 28963 7395
rect 30282 7392 30288 7404
rect 28951 7364 30288 7392
rect 28951 7361 28963 7364
rect 28905 7355 28963 7361
rect 30282 7352 30288 7364
rect 30340 7352 30346 7404
rect 32122 7392 32128 7404
rect 32083 7364 32128 7392
rect 32122 7352 32128 7364
rect 32180 7352 32186 7404
rect 33410 7352 33416 7404
rect 33468 7392 33474 7404
rect 33962 7392 33968 7404
rect 33468 7364 33968 7392
rect 33468 7352 33474 7364
rect 33962 7352 33968 7364
rect 34020 7392 34026 7404
rect 34425 7395 34483 7401
rect 34020 7364 34284 7392
rect 34020 7352 34026 7364
rect 18616 7296 22094 7324
rect 18233 7287 18291 7293
rect 9769 7259 9827 7265
rect 9769 7225 9781 7259
rect 9815 7256 9827 7259
rect 17954 7256 17960 7268
rect 9815 7228 17960 7256
rect 9815 7225 9827 7228
rect 9769 7219 9827 7225
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 18248 7256 18276 7287
rect 23474 7284 23480 7336
rect 23532 7324 23538 7336
rect 24029 7327 24087 7333
rect 24029 7324 24041 7327
rect 23532 7296 24041 7324
rect 23532 7284 23538 7296
rect 24029 7293 24041 7296
rect 24075 7293 24087 7327
rect 24029 7287 24087 7293
rect 30929 7327 30987 7333
rect 30929 7293 30941 7327
rect 30975 7324 30987 7327
rect 31478 7324 31484 7336
rect 30975 7296 31484 7324
rect 30975 7293 30987 7296
rect 30929 7287 30987 7293
rect 31478 7284 31484 7296
rect 31536 7284 31542 7336
rect 34149 7327 34207 7333
rect 34149 7324 34161 7327
rect 33980 7296 34161 7324
rect 20714 7256 20720 7268
rect 18248 7228 20720 7256
rect 20714 7216 20720 7228
rect 20772 7216 20778 7268
rect 10965 7191 11023 7197
rect 10965 7157 10977 7191
rect 11011 7188 11023 7191
rect 11514 7188 11520 7200
rect 11011 7160 11520 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 11514 7148 11520 7160
rect 11572 7148 11578 7200
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 12989 7191 13047 7197
rect 12989 7188 13001 7191
rect 12676 7160 13001 7188
rect 12676 7148 12682 7160
rect 12989 7157 13001 7160
rect 13035 7157 13047 7191
rect 12989 7151 13047 7157
rect 13633 7191 13691 7197
rect 13633 7157 13645 7191
rect 13679 7188 13691 7191
rect 14090 7188 14096 7200
rect 13679 7160 14096 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 17494 7148 17500 7200
rect 17552 7188 17558 7200
rect 25409 7191 25467 7197
rect 25409 7188 25421 7191
rect 17552 7160 25421 7188
rect 17552 7148 17558 7160
rect 25409 7157 25421 7160
rect 25455 7157 25467 7191
rect 25409 7151 25467 7157
rect 31294 7148 31300 7200
rect 31352 7188 31358 7200
rect 31389 7191 31447 7197
rect 31389 7188 31401 7191
rect 31352 7160 31401 7188
rect 31352 7148 31358 7160
rect 31389 7157 31401 7160
rect 31435 7157 31447 7191
rect 32306 7188 32312 7200
rect 32267 7160 32312 7188
rect 31389 7151 31447 7157
rect 32306 7148 32312 7160
rect 32364 7148 32370 7200
rect 32766 7188 32772 7200
rect 32727 7160 32772 7188
rect 32766 7148 32772 7160
rect 32824 7148 32830 7200
rect 33597 7191 33655 7197
rect 33597 7157 33609 7191
rect 33643 7188 33655 7191
rect 33980 7188 34008 7296
rect 34149 7293 34161 7296
rect 34195 7293 34207 7327
rect 34256 7324 34284 7364
rect 34425 7361 34437 7395
rect 34471 7392 34483 7395
rect 35986 7392 35992 7404
rect 34471 7364 35992 7392
rect 34471 7361 34483 7364
rect 34425 7355 34483 7361
rect 35986 7352 35992 7364
rect 36044 7352 36050 7404
rect 37829 7327 37887 7333
rect 37829 7324 37841 7327
rect 34256 7296 37841 7324
rect 34149 7287 34207 7293
rect 37829 7293 37841 7296
rect 37875 7293 37887 7327
rect 37829 7287 37887 7293
rect 34054 7216 34060 7268
rect 34112 7256 34118 7268
rect 35805 7259 35863 7265
rect 35805 7256 35817 7259
rect 34112 7228 35817 7256
rect 34112 7216 34118 7228
rect 35805 7225 35817 7228
rect 35851 7225 35863 7259
rect 35805 7219 35863 7225
rect 35894 7216 35900 7268
rect 35952 7256 35958 7268
rect 37277 7259 37335 7265
rect 37277 7256 37289 7259
rect 35952 7228 37289 7256
rect 35952 7216 35958 7228
rect 37277 7225 37289 7228
rect 37323 7225 37335 7259
rect 37277 7219 37335 7225
rect 35342 7188 35348 7200
rect 33643 7160 35348 7188
rect 33643 7157 33655 7160
rect 33597 7151 33655 7157
rect 35342 7148 35348 7160
rect 35400 7148 35406 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 15930 6984 15936 6996
rect 15891 6956 15936 6984
rect 15930 6944 15936 6956
rect 15988 6984 15994 6996
rect 15988 6956 16436 6984
rect 15988 6944 15994 6956
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12492 6820 12541 6848
rect 12492 6808 12498 6820
rect 12529 6817 12541 6820
rect 12575 6848 12587 6851
rect 12575 6820 13860 6848
rect 12575 6817 12587 6820
rect 12529 6811 12587 6817
rect 11514 6780 11520 6792
rect 11475 6752 11520 6780
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 12342 6740 12348 6792
rect 12400 6780 12406 6792
rect 13081 6783 13139 6789
rect 13081 6780 13093 6783
rect 12400 6752 13093 6780
rect 12400 6740 12406 6752
rect 13081 6749 13093 6752
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 12618 6672 12624 6724
rect 12676 6712 12682 6724
rect 13357 6715 13415 6721
rect 13357 6712 13369 6715
rect 12676 6684 13369 6712
rect 12676 6672 12682 6684
rect 13357 6681 13369 6684
rect 13403 6681 13415 6715
rect 13832 6712 13860 6820
rect 14090 6808 14096 6860
rect 14148 6848 14154 6860
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 14148 6820 14289 6848
rect 14148 6808 14154 6820
rect 14277 6817 14289 6820
rect 14323 6817 14335 6851
rect 14458 6848 14464 6860
rect 14419 6820 14464 6848
rect 14277 6811 14335 6817
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 15381 6851 15439 6857
rect 15381 6817 15393 6851
rect 15427 6848 15439 6851
rect 15562 6848 15568 6860
rect 15427 6820 15568 6848
rect 15427 6817 15439 6820
rect 15381 6811 15439 6817
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 16408 6857 16436 6956
rect 16942 6944 16948 6996
rect 17000 6984 17006 6996
rect 17865 6987 17923 6993
rect 17865 6984 17877 6987
rect 17000 6956 17877 6984
rect 17000 6944 17006 6956
rect 17865 6953 17877 6956
rect 17911 6953 17923 6987
rect 19242 6984 19248 6996
rect 19203 6956 19248 6984
rect 17865 6947 17923 6953
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 19334 6876 19340 6928
rect 19392 6916 19398 6928
rect 31665 6919 31723 6925
rect 19392 6888 19932 6916
rect 19392 6876 19398 6888
rect 16393 6851 16451 6857
rect 16393 6817 16405 6851
rect 16439 6817 16451 6851
rect 16393 6811 16451 6817
rect 18693 6851 18751 6857
rect 18693 6817 18705 6851
rect 18739 6848 18751 6851
rect 19150 6848 19156 6860
rect 18739 6820 19156 6848
rect 18739 6817 18751 6820
rect 18693 6811 18751 6817
rect 19150 6808 19156 6820
rect 19208 6848 19214 6860
rect 19797 6851 19855 6857
rect 19797 6848 19809 6851
rect 19208 6820 19809 6848
rect 19208 6808 19214 6820
rect 19797 6817 19809 6820
rect 19843 6817 19855 6851
rect 19904 6848 19932 6888
rect 31665 6885 31677 6919
rect 31711 6885 31723 6919
rect 31665 6879 31723 6885
rect 21726 6848 21732 6860
rect 19904 6820 21732 6848
rect 19797 6811 19855 6817
rect 21726 6808 21732 6820
rect 21784 6808 21790 6860
rect 30558 6848 30564 6860
rect 29932 6820 30564 6848
rect 13906 6740 13912 6792
rect 13964 6780 13970 6792
rect 14369 6783 14427 6789
rect 14369 6780 14381 6783
rect 13964 6752 14381 6780
rect 13964 6740 13970 6752
rect 14369 6749 14381 6752
rect 14415 6749 14427 6783
rect 14369 6743 14427 6749
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 15580 6780 15608 6808
rect 16577 6783 16635 6789
rect 16577 6780 16589 6783
rect 15580 6752 16589 6780
rect 14553 6743 14611 6749
rect 16577 6749 16589 6752
rect 16623 6749 16635 6783
rect 16577 6743 16635 6749
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6780 16819 6783
rect 17221 6783 17279 6789
rect 17221 6780 17233 6783
rect 16807 6752 17233 6780
rect 16807 6749 16819 6752
rect 16761 6743 16819 6749
rect 17221 6749 17233 6752
rect 17267 6749 17279 6783
rect 17221 6743 17279 6749
rect 14568 6712 14596 6743
rect 20070 6740 20076 6792
rect 20128 6780 20134 6792
rect 20441 6783 20499 6789
rect 20441 6780 20453 6783
rect 20128 6752 20453 6780
rect 20128 6740 20134 6752
rect 20441 6749 20453 6752
rect 20487 6749 20499 6783
rect 20441 6743 20499 6749
rect 22186 6740 22192 6792
rect 22244 6780 22250 6792
rect 23017 6783 23075 6789
rect 22244 6752 22876 6780
rect 22244 6740 22250 6752
rect 16390 6712 16396 6724
rect 13832 6684 16396 6712
rect 13357 6675 13415 6681
rect 16390 6672 16396 6684
rect 16448 6672 16454 6724
rect 19334 6672 19340 6724
rect 19392 6712 19398 6724
rect 19518 6712 19524 6724
rect 19392 6684 19524 6712
rect 19392 6672 19398 6684
rect 19518 6672 19524 6684
rect 19576 6672 19582 6724
rect 22278 6712 22284 6724
rect 20640 6684 22284 6712
rect 11054 6644 11060 6656
rect 11015 6616 11060 6644
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11698 6644 11704 6656
rect 11659 6616 11704 6644
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 14090 6644 14096 6656
rect 14051 6616 14096 6644
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 17402 6644 17408 6656
rect 17363 6616 17408 6644
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 18966 6604 18972 6656
rect 19024 6644 19030 6656
rect 19613 6647 19671 6653
rect 19613 6644 19625 6647
rect 19024 6616 19625 6644
rect 19024 6604 19030 6616
rect 19613 6613 19625 6616
rect 19659 6613 19671 6647
rect 19613 6607 19671 6613
rect 19705 6647 19763 6653
rect 19705 6613 19717 6647
rect 19751 6644 19763 6647
rect 20162 6644 20168 6656
rect 19751 6616 20168 6644
rect 19751 6613 19763 6616
rect 19705 6607 19763 6613
rect 20162 6604 20168 6616
rect 20220 6604 20226 6656
rect 20640 6653 20668 6684
rect 22278 6672 22284 6684
rect 22336 6672 22342 6724
rect 22750 6715 22808 6721
rect 22750 6712 22762 6715
rect 22388 6684 22762 6712
rect 20625 6647 20683 6653
rect 20625 6613 20637 6647
rect 20671 6613 20683 6647
rect 21634 6644 21640 6656
rect 21595 6616 21640 6644
rect 20625 6607 20683 6613
rect 21634 6604 21640 6616
rect 21692 6604 21698 6656
rect 21726 6604 21732 6656
rect 21784 6644 21790 6656
rect 22388 6644 22416 6684
rect 22750 6681 22762 6684
rect 22796 6681 22808 6715
rect 22750 6675 22808 6681
rect 21784 6616 22416 6644
rect 22848 6644 22876 6752
rect 23017 6749 23029 6783
rect 23063 6780 23075 6783
rect 23474 6780 23480 6792
rect 23063 6752 23480 6780
rect 23063 6749 23075 6752
rect 23017 6743 23075 6749
rect 23474 6740 23480 6752
rect 23532 6740 23538 6792
rect 23566 6740 23572 6792
rect 23624 6780 23630 6792
rect 26890 6783 26948 6789
rect 26890 6780 26902 6783
rect 23624 6752 26902 6780
rect 23624 6740 23630 6752
rect 26890 6749 26902 6752
rect 26936 6749 26948 6783
rect 26890 6743 26948 6749
rect 27157 6783 27215 6789
rect 27157 6749 27169 6783
rect 27203 6780 27215 6783
rect 27614 6780 27620 6792
rect 27203 6752 27620 6780
rect 27203 6749 27215 6752
rect 27157 6743 27215 6749
rect 27614 6740 27620 6752
rect 27672 6780 27678 6792
rect 28350 6780 28356 6792
rect 27672 6752 28356 6780
rect 27672 6740 27678 6752
rect 28350 6740 28356 6752
rect 28408 6740 28414 6792
rect 24762 6672 24768 6724
rect 24820 6712 24826 6724
rect 29932 6721 29960 6820
rect 30558 6808 30564 6820
rect 30616 6808 30622 6860
rect 30742 6848 30748 6860
rect 30703 6820 30748 6848
rect 30742 6808 30748 6820
rect 30800 6848 30806 6860
rect 31680 6848 31708 6879
rect 30800 6820 31708 6848
rect 30800 6808 30806 6820
rect 34330 6808 34336 6860
rect 34388 6848 34394 6860
rect 35161 6851 35219 6857
rect 35161 6848 35173 6851
rect 34388 6820 35173 6848
rect 34388 6808 34394 6820
rect 35161 6817 35173 6820
rect 35207 6817 35219 6851
rect 35342 6848 35348 6860
rect 35303 6820 35348 6848
rect 35161 6811 35219 6817
rect 35342 6808 35348 6820
rect 35400 6808 35406 6860
rect 36170 6848 36176 6860
rect 36131 6820 36176 6848
rect 36170 6808 36176 6820
rect 36228 6808 36234 6860
rect 31478 6740 31484 6792
rect 31536 6780 31542 6792
rect 33045 6783 33103 6789
rect 33045 6780 33057 6783
rect 31536 6752 33057 6780
rect 31536 6740 31542 6752
rect 33045 6749 33057 6752
rect 33091 6749 33103 6783
rect 33962 6780 33968 6792
rect 33923 6752 33968 6780
rect 33045 6743 33103 6749
rect 33962 6740 33968 6752
rect 34020 6740 34026 6792
rect 35069 6783 35127 6789
rect 35069 6749 35081 6783
rect 35115 6780 35127 6783
rect 37182 6780 37188 6792
rect 35115 6752 37188 6780
rect 35115 6749 35127 6752
rect 35069 6743 35127 6749
rect 37182 6740 37188 6752
rect 37240 6740 37246 6792
rect 29917 6715 29975 6721
rect 29917 6712 29929 6715
rect 24820 6684 29929 6712
rect 24820 6672 24826 6684
rect 29917 6681 29929 6684
rect 29963 6681 29975 6715
rect 29917 6675 29975 6681
rect 31220 6684 31754 6712
rect 25777 6647 25835 6653
rect 25777 6644 25789 6647
rect 22848 6616 25789 6644
rect 21784 6604 21790 6616
rect 25777 6613 25789 6616
rect 25823 6613 25835 6647
rect 25777 6607 25835 6613
rect 30834 6604 30840 6656
rect 30892 6644 30898 6656
rect 31220 6653 31248 6684
rect 31205 6647 31263 6653
rect 30892 6616 30937 6644
rect 30892 6604 30898 6616
rect 31205 6613 31217 6647
rect 31251 6613 31263 6647
rect 31726 6644 31754 6684
rect 32306 6672 32312 6724
rect 32364 6712 32370 6724
rect 32778 6715 32836 6721
rect 32778 6712 32790 6715
rect 32364 6684 32790 6712
rect 32364 6672 32370 6684
rect 32778 6681 32790 6684
rect 32824 6681 32836 6715
rect 36418 6715 36476 6721
rect 36418 6712 36430 6715
rect 32778 6675 32836 6681
rect 34164 6684 36430 6712
rect 32122 6644 32128 6656
rect 31726 6616 32128 6644
rect 31205 6607 31263 6613
rect 32122 6604 32128 6616
rect 32180 6604 32186 6656
rect 34164 6653 34192 6684
rect 36418 6681 36430 6684
rect 36464 6681 36476 6715
rect 38013 6715 38071 6721
rect 38013 6712 38025 6715
rect 36418 6675 36476 6681
rect 36556 6684 38025 6712
rect 34149 6647 34207 6653
rect 34149 6613 34161 6647
rect 34195 6613 34207 6647
rect 34149 6607 34207 6613
rect 34422 6604 34428 6656
rect 34480 6644 34486 6656
rect 34701 6647 34759 6653
rect 34701 6644 34713 6647
rect 34480 6616 34713 6644
rect 34480 6604 34486 6616
rect 34701 6613 34713 6616
rect 34747 6613 34759 6647
rect 34701 6607 34759 6613
rect 36078 6604 36084 6656
rect 36136 6644 36142 6656
rect 36556 6644 36584 6684
rect 38013 6681 38025 6684
rect 38059 6681 38071 6715
rect 38013 6675 38071 6681
rect 37550 6644 37556 6656
rect 36136 6616 36584 6644
rect 37511 6616 37556 6644
rect 36136 6604 36142 6616
rect 37550 6604 37556 6616
rect 37608 6604 37614 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 9953 6443 10011 6449
rect 9953 6440 9965 6443
rect 9732 6412 9965 6440
rect 9732 6400 9738 6412
rect 9953 6409 9965 6412
rect 9999 6409 10011 6443
rect 11885 6443 11943 6449
rect 11885 6440 11897 6443
rect 9953 6403 10011 6409
rect 10152 6412 11897 6440
rect 8386 6332 8392 6384
rect 8444 6372 8450 6384
rect 10152 6372 10180 6412
rect 11885 6409 11897 6412
rect 11931 6409 11943 6443
rect 11885 6403 11943 6409
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 12253 6443 12311 6449
rect 12253 6440 12265 6443
rect 12216 6412 12265 6440
rect 12216 6400 12222 6412
rect 12253 6409 12265 6412
rect 12299 6409 12311 6443
rect 13906 6440 13912 6452
rect 13867 6412 13912 6440
rect 12253 6403 12311 6409
rect 13906 6400 13912 6412
rect 13964 6400 13970 6452
rect 18966 6440 18972 6452
rect 16592 6412 18972 6440
rect 8444 6344 10180 6372
rect 8444 6332 8450 6344
rect 10410 6332 10416 6384
rect 10468 6372 10474 6384
rect 10505 6375 10563 6381
rect 10505 6372 10517 6375
rect 10468 6344 10517 6372
rect 10468 6332 10474 6344
rect 10505 6341 10517 6344
rect 10551 6341 10563 6375
rect 10505 6335 10563 6341
rect 11793 6375 11851 6381
rect 11793 6341 11805 6375
rect 11839 6372 11851 6375
rect 12066 6372 12072 6384
rect 11839 6344 12072 6372
rect 11839 6341 11851 6344
rect 11793 6335 11851 6341
rect 10520 6236 10548 6335
rect 12066 6332 12072 6344
rect 12124 6372 12130 6384
rect 12526 6372 12532 6384
rect 12124 6344 12532 6372
rect 12124 6332 12130 6344
rect 12526 6332 12532 6344
rect 12584 6372 12590 6384
rect 13354 6372 13360 6384
rect 12584 6344 13360 6372
rect 12584 6332 12590 6344
rect 13354 6332 13360 6344
rect 13412 6332 13418 6384
rect 14737 6375 14795 6381
rect 14737 6372 14749 6375
rect 13648 6344 14749 6372
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6304 10931 6307
rect 11698 6304 11704 6316
rect 10919 6276 11704 6304
rect 10919 6273 10931 6276
rect 10873 6267 10931 6273
rect 11698 6264 11704 6276
rect 11756 6304 11762 6316
rect 11756 6276 11836 6304
rect 11756 6264 11762 6276
rect 11609 6239 11667 6245
rect 11609 6236 11621 6239
rect 10520 6208 11621 6236
rect 11609 6205 11621 6208
rect 11655 6205 11667 6239
rect 11808 6236 11836 6276
rect 12618 6264 12624 6316
rect 12676 6304 12682 6316
rect 12713 6307 12771 6313
rect 12713 6304 12725 6307
rect 12676 6276 12725 6304
rect 12676 6264 12682 6276
rect 12713 6273 12725 6276
rect 12759 6273 12771 6307
rect 12713 6267 12771 6273
rect 12894 6264 12900 6316
rect 12952 6304 12958 6316
rect 13170 6304 13176 6316
rect 12952 6276 13176 6304
rect 12952 6264 12958 6276
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 13538 6304 13544 6316
rect 13499 6276 13544 6304
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 12342 6236 12348 6248
rect 11808 6208 12348 6236
rect 11609 6199 11667 6205
rect 12342 6196 12348 6208
rect 12400 6236 12406 6248
rect 13648 6236 13676 6344
rect 14737 6341 14749 6344
rect 14783 6341 14795 6375
rect 14737 6335 14795 6341
rect 15105 6375 15163 6381
rect 15105 6341 15117 6375
rect 15151 6372 15163 6375
rect 16482 6372 16488 6384
rect 15151 6344 16488 6372
rect 15151 6341 15163 6344
rect 15105 6335 15163 6341
rect 13722 6264 13728 6316
rect 13780 6304 13786 6316
rect 14752 6304 14780 6335
rect 16482 6332 16488 6344
rect 16540 6332 16546 6384
rect 15749 6307 15807 6313
rect 15749 6304 15761 6307
rect 13780 6276 13873 6304
rect 14752 6276 15761 6304
rect 13780 6264 13786 6276
rect 15749 6273 15761 6276
rect 15795 6273 15807 6307
rect 16114 6304 16120 6316
rect 16027 6276 16120 6304
rect 15749 6267 15807 6273
rect 12400 6208 13676 6236
rect 12400 6196 12406 6208
rect 13740 6168 13768 6264
rect 15764 6236 15792 6267
rect 16114 6264 16120 6276
rect 16172 6304 16178 6316
rect 16592 6304 16620 6412
rect 18966 6400 18972 6412
rect 19024 6400 19030 6452
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 19392 6412 19441 6440
rect 19392 6400 19398 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 20162 6440 20168 6452
rect 20075 6412 20168 6440
rect 19429 6403 19487 6409
rect 20162 6400 20168 6412
rect 20220 6440 20226 6452
rect 22278 6440 22284 6452
rect 20220 6412 22284 6440
rect 20220 6400 20226 6412
rect 22278 6400 22284 6412
rect 22336 6400 22342 6452
rect 22370 6400 22376 6452
rect 22428 6440 22434 6452
rect 28445 6443 28503 6449
rect 28445 6440 28457 6443
rect 22428 6412 28457 6440
rect 22428 6400 22434 6412
rect 28445 6409 28457 6412
rect 28491 6409 28503 6443
rect 28445 6403 28503 6409
rect 28810 6400 28816 6452
rect 28868 6440 28874 6452
rect 30282 6440 30288 6452
rect 28868 6412 30144 6440
rect 30243 6412 30288 6440
rect 28868 6400 28874 6412
rect 18138 6372 18144 6384
rect 16776 6344 18144 6372
rect 16776 6313 16804 6344
rect 18138 6332 18144 6344
rect 18196 6332 18202 6384
rect 18325 6375 18383 6381
rect 18325 6341 18337 6375
rect 18371 6372 18383 6375
rect 24734 6375 24792 6381
rect 24734 6372 24746 6375
rect 18371 6344 24746 6372
rect 18371 6341 18383 6344
rect 18325 6335 18383 6341
rect 24734 6341 24746 6344
rect 24780 6341 24792 6375
rect 24734 6335 24792 6341
rect 28350 6332 28356 6384
rect 28408 6372 28414 6384
rect 30116 6372 30144 6412
rect 30282 6400 30288 6412
rect 30340 6400 30346 6452
rect 30745 6443 30803 6449
rect 30745 6440 30757 6443
rect 30484 6412 30757 6440
rect 30484 6372 30512 6412
rect 30745 6409 30757 6412
rect 30791 6440 30803 6443
rect 31386 6440 31392 6452
rect 30791 6412 31392 6440
rect 30791 6409 30803 6412
rect 30745 6403 30803 6409
rect 31386 6400 31392 6412
rect 31444 6400 31450 6452
rect 32401 6443 32459 6449
rect 32401 6409 32413 6443
rect 32447 6440 32459 6443
rect 32490 6440 32496 6452
rect 32447 6412 32496 6440
rect 32447 6409 32459 6412
rect 32401 6403 32459 6409
rect 32490 6400 32496 6412
rect 32548 6400 32554 6452
rect 32861 6443 32919 6449
rect 32861 6409 32873 6443
rect 32907 6440 32919 6443
rect 33962 6440 33968 6452
rect 32907 6412 33968 6440
rect 32907 6409 32919 6412
rect 32861 6403 32919 6409
rect 33962 6400 33968 6412
rect 34020 6400 34026 6452
rect 34330 6400 34336 6452
rect 34388 6440 34394 6452
rect 35805 6443 35863 6449
rect 35805 6440 35817 6443
rect 34388 6412 35817 6440
rect 34388 6400 34394 6412
rect 35805 6409 35817 6412
rect 35851 6409 35863 6443
rect 35805 6403 35863 6409
rect 28408 6344 29868 6372
rect 30116 6344 30512 6372
rect 28408 6332 28414 6344
rect 16172 6276 16620 6304
rect 16761 6307 16819 6313
rect 16172 6264 16178 6276
rect 16761 6273 16773 6307
rect 16807 6273 16819 6307
rect 16761 6267 16819 6273
rect 16776 6236 16804 6267
rect 17034 6264 17040 6316
rect 17092 6304 17098 6316
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 17092 6276 18245 6304
rect 17092 6264 17098 6276
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18417 6307 18475 6313
rect 18417 6304 18429 6307
rect 18233 6267 18291 6273
rect 18340 6276 18429 6304
rect 15764 6208 16804 6236
rect 16850 6196 16856 6248
rect 16908 6236 16914 6248
rect 16945 6239 17003 6245
rect 16945 6236 16957 6239
rect 16908 6208 16957 6236
rect 16908 6196 16914 6208
rect 16945 6205 16957 6208
rect 16991 6236 17003 6239
rect 17770 6236 17776 6248
rect 16991 6208 17776 6236
rect 16991 6205 17003 6208
rect 16945 6199 17003 6205
rect 17770 6196 17776 6208
rect 17828 6196 17834 6248
rect 17310 6168 17316 6180
rect 13740 6140 17316 6168
rect 17310 6128 17316 6140
rect 17368 6128 17374 6180
rect 18340 6168 18368 6276
rect 18417 6273 18429 6276
rect 18463 6273 18475 6307
rect 18417 6267 18475 6273
rect 18598 6264 18604 6316
rect 18656 6304 18662 6316
rect 22934 6307 22992 6313
rect 22934 6304 22946 6307
rect 18656 6276 22946 6304
rect 18656 6264 18662 6276
rect 22934 6273 22946 6276
rect 22980 6273 22992 6307
rect 22934 6267 22992 6273
rect 28994 6264 29000 6316
rect 29052 6304 29058 6316
rect 29840 6313 29868 6344
rect 30558 6332 30564 6384
rect 30616 6372 30622 6384
rect 31481 6375 31539 6381
rect 31481 6372 31493 6375
rect 30616 6344 31493 6372
rect 30616 6332 30622 6344
rect 29558 6307 29616 6313
rect 29558 6304 29570 6307
rect 29052 6276 29570 6304
rect 29052 6264 29058 6276
rect 29558 6273 29570 6276
rect 29604 6273 29616 6307
rect 29558 6267 29616 6273
rect 29825 6307 29883 6313
rect 29825 6273 29837 6307
rect 29871 6273 29883 6307
rect 30650 6304 30656 6316
rect 30611 6276 30656 6304
rect 29825 6267 29883 6273
rect 30650 6264 30656 6276
rect 30708 6264 30714 6316
rect 23201 6239 23259 6245
rect 23201 6205 23213 6239
rect 23247 6236 23259 6239
rect 23474 6236 23480 6248
rect 23247 6208 23480 6236
rect 23247 6205 23259 6208
rect 23201 6199 23259 6205
rect 23474 6196 23480 6208
rect 23532 6236 23538 6248
rect 30852 6245 30880 6344
rect 31481 6341 31493 6344
rect 31527 6372 31539 6375
rect 33226 6372 33232 6384
rect 31527 6344 31754 6372
rect 31527 6341 31539 6344
rect 31481 6335 31539 6341
rect 24489 6239 24547 6245
rect 24489 6236 24501 6239
rect 23532 6208 24501 6236
rect 23532 6196 23538 6208
rect 24489 6205 24501 6208
rect 24535 6205 24547 6239
rect 24489 6199 24547 6205
rect 30837 6239 30895 6245
rect 30837 6205 30849 6239
rect 30883 6205 30895 6239
rect 31726 6236 31754 6344
rect 32324 6344 33232 6372
rect 32030 6236 32036 6248
rect 31726 6208 32036 6236
rect 30837 6199 30895 6205
rect 32030 6196 32036 6208
rect 32088 6236 32094 6248
rect 32324 6245 32352 6344
rect 33226 6332 33232 6344
rect 33284 6332 33290 6384
rect 32493 6307 32551 6313
rect 32493 6273 32505 6307
rect 32539 6304 32551 6307
rect 33962 6304 33968 6316
rect 32539 6276 33968 6304
rect 32539 6273 32551 6276
rect 32493 6267 32551 6273
rect 33962 6264 33968 6276
rect 34020 6264 34026 6316
rect 34609 6307 34667 6313
rect 34609 6273 34621 6307
rect 34655 6304 34667 6307
rect 34698 6304 34704 6316
rect 34655 6276 34704 6304
rect 34655 6273 34667 6276
rect 34609 6267 34667 6273
rect 34698 6264 34704 6276
rect 34756 6264 34762 6316
rect 37645 6307 37703 6313
rect 37645 6273 37657 6307
rect 37691 6273 37703 6307
rect 37645 6267 37703 6273
rect 32309 6239 32367 6245
rect 32309 6236 32321 6239
rect 32088 6208 32321 6236
rect 32088 6196 32094 6208
rect 32309 6205 32321 6208
rect 32355 6205 32367 6239
rect 32309 6199 32367 6205
rect 33686 6196 33692 6248
rect 33744 6236 33750 6248
rect 37660 6236 37688 6267
rect 33744 6208 37688 6236
rect 33744 6196 33750 6208
rect 20254 6168 20260 6180
rect 17696 6140 20260 6168
rect 12526 6060 12532 6112
rect 12584 6100 12590 6112
rect 12713 6103 12771 6109
rect 12713 6100 12725 6103
rect 12584 6072 12725 6100
rect 12584 6060 12590 6072
rect 12713 6069 12725 6072
rect 12759 6069 12771 6103
rect 15562 6100 15568 6112
rect 15523 6072 15568 6100
rect 12713 6063 12771 6069
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 15746 6100 15752 6112
rect 15707 6072 15752 6100
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 17696 6109 17724 6140
rect 20254 6128 20260 6140
rect 20312 6128 20318 6180
rect 20438 6128 20444 6180
rect 20496 6168 20502 6180
rect 21085 6171 21143 6177
rect 21085 6168 21097 6171
rect 20496 6140 21097 6168
rect 20496 6128 20502 6140
rect 21085 6137 21097 6140
rect 21131 6168 21143 6171
rect 21450 6168 21456 6180
rect 21131 6140 21456 6168
rect 21131 6137 21143 6140
rect 21085 6131 21143 6137
rect 21450 6128 21456 6140
rect 21508 6128 21514 6180
rect 21560 6140 22094 6168
rect 17681 6103 17739 6109
rect 17681 6100 17693 6103
rect 16448 6072 17693 6100
rect 16448 6060 16454 6072
rect 17681 6069 17693 6072
rect 17727 6069 17739 6103
rect 17681 6063 17739 6069
rect 17770 6060 17776 6112
rect 17828 6100 17834 6112
rect 21560 6100 21588 6140
rect 21818 6100 21824 6112
rect 17828 6072 21588 6100
rect 21779 6072 21824 6100
rect 17828 6060 17834 6072
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 22066 6100 22094 6140
rect 32950 6128 32956 6180
rect 33008 6168 33014 6180
rect 33873 6171 33931 6177
rect 33873 6168 33885 6171
rect 33008 6140 33885 6168
rect 33008 6128 33014 6140
rect 33873 6137 33885 6140
rect 33919 6137 33931 6171
rect 37550 6168 37556 6180
rect 33873 6131 33931 6137
rect 34624 6140 37556 6168
rect 24762 6100 24768 6112
rect 22066 6072 24768 6100
rect 24762 6060 24768 6072
rect 24820 6060 24826 6112
rect 24854 6060 24860 6112
rect 24912 6100 24918 6112
rect 25869 6103 25927 6109
rect 25869 6100 25881 6103
rect 24912 6072 25881 6100
rect 24912 6060 24918 6072
rect 25869 6069 25881 6072
rect 25915 6069 25927 6103
rect 25869 6063 25927 6069
rect 32490 6060 32496 6112
rect 32548 6100 32554 6112
rect 33321 6103 33379 6109
rect 33321 6100 33333 6103
rect 32548 6072 33333 6100
rect 32548 6060 32554 6072
rect 33321 6069 33333 6072
rect 33367 6100 33379 6103
rect 34624 6100 34652 6140
rect 37550 6128 37556 6140
rect 37608 6128 37614 6180
rect 34790 6100 34796 6112
rect 33367 6072 34652 6100
rect 34751 6072 34796 6100
rect 33367 6069 33379 6072
rect 33321 6063 33379 6069
rect 34790 6060 34796 6072
rect 34848 6060 34854 6112
rect 35342 6100 35348 6112
rect 35303 6072 35348 6100
rect 35342 6060 35348 6072
rect 35400 6100 35406 6112
rect 36357 6103 36415 6109
rect 36357 6100 36369 6103
rect 35400 6072 36369 6100
rect 35400 6060 35406 6072
rect 36357 6069 36369 6072
rect 36403 6069 36415 6103
rect 36357 6063 36415 6069
rect 36630 6060 36636 6112
rect 36688 6100 36694 6112
rect 37461 6103 37519 6109
rect 37461 6100 37473 6103
rect 36688 6072 37473 6100
rect 36688 6060 36694 6072
rect 37461 6069 37473 6072
rect 37507 6069 37519 6103
rect 37461 6063 37519 6069
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 9950 5896 9956 5908
rect 9911 5868 9956 5896
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 12066 5896 12072 5908
rect 12027 5868 12072 5896
rect 12066 5856 12072 5868
rect 12124 5856 12130 5908
rect 12894 5896 12900 5908
rect 12855 5868 12900 5896
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 15473 5899 15531 5905
rect 15473 5896 15485 5899
rect 13044 5868 15485 5896
rect 13044 5856 13050 5868
rect 15473 5865 15485 5868
rect 15519 5896 15531 5899
rect 16114 5896 16120 5908
rect 15519 5868 16120 5896
rect 15519 5865 15531 5868
rect 15473 5859 15531 5865
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 17313 5899 17371 5905
rect 17313 5865 17325 5899
rect 17359 5896 17371 5899
rect 19426 5896 19432 5908
rect 17359 5868 19432 5896
rect 17359 5865 17371 5868
rect 17313 5859 17371 5865
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 19996 5868 25820 5896
rect 11057 5831 11115 5837
rect 11057 5797 11069 5831
rect 11103 5828 11115 5831
rect 18598 5828 18604 5840
rect 11103 5800 18604 5828
rect 11103 5797 11115 5800
rect 11057 5791 11115 5797
rect 18598 5788 18604 5800
rect 18656 5788 18662 5840
rect 19334 5788 19340 5840
rect 19392 5828 19398 5840
rect 19996 5828 20024 5868
rect 20530 5828 20536 5840
rect 19392 5800 20024 5828
rect 20491 5800 20536 5828
rect 19392 5788 19398 5800
rect 20530 5788 20536 5800
rect 20588 5788 20594 5840
rect 22097 5831 22155 5837
rect 22097 5828 22109 5831
rect 20640 5800 22109 5828
rect 9401 5763 9459 5769
rect 9401 5729 9413 5763
rect 9447 5729 9459 5763
rect 9401 5723 9459 5729
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5760 9551 5763
rect 9674 5760 9680 5772
rect 9539 5732 9680 5760
rect 9539 5729 9551 5732
rect 9493 5723 9551 5729
rect 9416 5692 9444 5723
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 13170 5720 13176 5772
rect 13228 5760 13234 5772
rect 13357 5763 13415 5769
rect 13357 5760 13369 5763
rect 13228 5732 13369 5760
rect 13228 5720 13234 5732
rect 13357 5729 13369 5732
rect 13403 5760 13415 5763
rect 15746 5760 15752 5772
rect 13403 5732 15752 5760
rect 13403 5729 13415 5732
rect 13357 5723 13415 5729
rect 15746 5720 15752 5732
rect 15804 5760 15810 5772
rect 16025 5763 16083 5769
rect 16025 5760 16037 5763
rect 15804 5732 16037 5760
rect 15804 5720 15810 5732
rect 16025 5729 16037 5732
rect 16071 5729 16083 5763
rect 16025 5723 16083 5729
rect 16482 5720 16488 5772
rect 16540 5760 16546 5772
rect 16669 5763 16727 5769
rect 16669 5760 16681 5763
rect 16540 5732 16681 5760
rect 16540 5720 16546 5732
rect 16669 5729 16681 5732
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 17494 5720 17500 5772
rect 17552 5760 17558 5772
rect 18693 5763 18751 5769
rect 18693 5760 18705 5763
rect 17552 5732 18705 5760
rect 17552 5720 17558 5732
rect 18693 5729 18705 5732
rect 18739 5729 18751 5763
rect 18693 5723 18751 5729
rect 10410 5692 10416 5704
rect 9416 5664 10416 5692
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 10870 5692 10876 5704
rect 10831 5664 10876 5692
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5692 12679 5695
rect 12710 5692 12716 5704
rect 12667 5664 12716 5692
rect 12667 5661 12679 5664
rect 12621 5655 12679 5661
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 12897 5695 12955 5701
rect 12897 5661 12909 5695
rect 12943 5692 12955 5695
rect 14090 5692 14096 5704
rect 12943 5664 14096 5692
rect 12943 5661 12955 5664
rect 12897 5655 12955 5661
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 14921 5695 14979 5701
rect 14921 5661 14933 5695
rect 14967 5692 14979 5695
rect 16850 5692 16856 5704
rect 14967 5664 16856 5692
rect 14967 5661 14979 5664
rect 14921 5655 14979 5661
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 17310 5652 17316 5704
rect 17368 5692 17374 5704
rect 18141 5695 18199 5701
rect 18141 5692 18153 5695
rect 17368 5664 18153 5692
rect 17368 5652 17374 5664
rect 18141 5661 18153 5664
rect 18187 5692 18199 5695
rect 20640 5692 20668 5800
rect 22097 5797 22109 5800
rect 22143 5797 22155 5831
rect 25792 5828 25820 5868
rect 26142 5856 26148 5908
rect 26200 5896 26206 5908
rect 26881 5899 26939 5905
rect 26881 5896 26893 5899
rect 26200 5868 26893 5896
rect 26200 5856 26206 5868
rect 26881 5865 26893 5868
rect 26927 5865 26939 5899
rect 29549 5899 29607 5905
rect 29549 5896 29561 5899
rect 26881 5859 26939 5865
rect 26988 5868 29561 5896
rect 26988 5828 27016 5868
rect 29549 5865 29561 5868
rect 29595 5865 29607 5899
rect 31386 5896 31392 5908
rect 31347 5868 31392 5896
rect 29549 5859 29607 5865
rect 31386 5856 31392 5868
rect 31444 5896 31450 5908
rect 33134 5896 33140 5908
rect 31444 5868 33140 5896
rect 31444 5856 31450 5868
rect 33134 5856 33140 5868
rect 33192 5856 33198 5908
rect 33226 5856 33232 5908
rect 33284 5896 33290 5908
rect 33597 5899 33655 5905
rect 33597 5896 33609 5899
rect 33284 5868 33609 5896
rect 33284 5856 33290 5868
rect 33597 5865 33609 5868
rect 33643 5865 33655 5899
rect 34698 5896 34704 5908
rect 34659 5868 34704 5896
rect 33597 5859 33655 5865
rect 34698 5856 34704 5868
rect 34756 5856 34762 5908
rect 35986 5896 35992 5908
rect 35947 5868 35992 5896
rect 35986 5856 35992 5868
rect 36044 5856 36050 5908
rect 37366 5896 37372 5908
rect 36096 5868 37372 5896
rect 25792 5800 27016 5828
rect 28997 5831 29055 5837
rect 22097 5791 22155 5797
rect 28997 5797 29009 5831
rect 29043 5828 29055 5831
rect 29178 5828 29184 5840
rect 29043 5800 29184 5828
rect 29043 5797 29055 5800
rect 28997 5791 29055 5797
rect 29178 5788 29184 5800
rect 29236 5788 29242 5840
rect 32030 5828 32036 5840
rect 31991 5800 32036 5828
rect 32030 5788 32036 5800
rect 32088 5788 32094 5840
rect 36096 5828 36124 5868
rect 37366 5856 37372 5868
rect 37424 5896 37430 5908
rect 38105 5899 38163 5905
rect 38105 5896 38117 5899
rect 37424 5868 38117 5896
rect 37424 5856 37430 5868
rect 38105 5865 38117 5868
rect 38151 5865 38163 5899
rect 38105 5859 38163 5865
rect 35176 5800 36124 5828
rect 35176 5769 35204 5800
rect 36170 5788 36176 5840
rect 36228 5828 36234 5840
rect 36228 5800 36768 5828
rect 36228 5788 36234 5800
rect 21361 5763 21419 5769
rect 21361 5760 21373 5763
rect 20824 5732 21373 5760
rect 20824 5701 20852 5732
rect 21361 5729 21373 5732
rect 21407 5729 21419 5763
rect 21361 5723 21419 5729
rect 35161 5763 35219 5769
rect 35161 5729 35173 5763
rect 35207 5729 35219 5763
rect 35342 5760 35348 5772
rect 35303 5732 35348 5760
rect 35161 5723 35219 5729
rect 35342 5720 35348 5732
rect 35400 5720 35406 5772
rect 36740 5769 36768 5800
rect 36725 5763 36783 5769
rect 36725 5729 36737 5763
rect 36771 5729 36783 5763
rect 36725 5723 36783 5729
rect 18187 5664 20668 5692
rect 20809 5695 20867 5701
rect 18187 5661 18199 5664
rect 18141 5655 18199 5661
rect 20809 5661 20821 5695
rect 20855 5661 20867 5695
rect 21266 5692 21272 5704
rect 21227 5664 21272 5692
rect 20809 5655 20867 5661
rect 21266 5652 21272 5664
rect 21324 5652 21330 5704
rect 21450 5692 21456 5704
rect 21411 5664 21456 5692
rect 21450 5652 21456 5664
rect 21508 5652 21514 5704
rect 22646 5652 22652 5704
rect 22704 5692 22710 5704
rect 23210 5695 23268 5701
rect 23210 5692 23222 5695
rect 22704 5664 23222 5692
rect 22704 5652 22710 5664
rect 23210 5661 23222 5664
rect 23256 5661 23268 5695
rect 23474 5692 23480 5704
rect 23435 5664 23480 5692
rect 23210 5655 23268 5661
rect 23474 5652 23480 5664
rect 23532 5652 23538 5704
rect 27614 5652 27620 5704
rect 27672 5692 27678 5704
rect 27994 5695 28052 5701
rect 27994 5692 28006 5695
rect 27672 5664 28006 5692
rect 27672 5652 27678 5664
rect 27994 5661 28006 5664
rect 28040 5661 28052 5695
rect 27994 5655 28052 5661
rect 28261 5695 28319 5701
rect 28261 5661 28273 5695
rect 28307 5692 28319 5695
rect 28350 5692 28356 5704
rect 28307 5664 28356 5692
rect 28307 5661 28319 5664
rect 28261 5655 28319 5661
rect 28350 5652 28356 5664
rect 28408 5652 28414 5704
rect 29638 5652 29644 5704
rect 29696 5692 29702 5704
rect 30929 5695 30987 5701
rect 29696 5664 30788 5692
rect 29696 5652 29702 5664
rect 8478 5584 8484 5636
rect 8536 5624 8542 5636
rect 9585 5627 9643 5633
rect 9585 5624 9597 5627
rect 8536 5596 9597 5624
rect 8536 5584 8542 5596
rect 9585 5593 9597 5596
rect 9631 5593 9643 5627
rect 9585 5587 9643 5593
rect 11609 5627 11667 5633
rect 11609 5593 11621 5627
rect 11655 5624 11667 5627
rect 13998 5624 14004 5636
rect 11655 5596 14004 5624
rect 11655 5593 11667 5596
rect 11609 5587 11667 5593
rect 13998 5584 14004 5596
rect 14056 5584 14062 5636
rect 14458 5584 14464 5636
rect 14516 5624 14522 5636
rect 16945 5627 17003 5633
rect 16945 5624 16957 5627
rect 14516 5596 16957 5624
rect 14516 5584 14522 5596
rect 16945 5593 16957 5596
rect 16991 5593 17003 5627
rect 17494 5624 17500 5636
rect 16945 5587 17003 5593
rect 17144 5596 17500 5624
rect 7929 5559 7987 5565
rect 7929 5525 7941 5559
rect 7975 5556 7987 5559
rect 8294 5556 8300 5568
rect 7975 5528 8300 5556
rect 7975 5525 7987 5528
rect 7929 5519 7987 5525
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 12526 5516 12532 5568
rect 12584 5556 12590 5568
rect 12713 5559 12771 5565
rect 12713 5556 12725 5559
rect 12584 5528 12725 5556
rect 12584 5516 12590 5528
rect 12713 5525 12725 5528
rect 12759 5525 12771 5559
rect 12713 5519 12771 5525
rect 14369 5559 14427 5565
rect 14369 5525 14381 5559
rect 14415 5556 14427 5559
rect 14734 5556 14740 5568
rect 14415 5528 14740 5556
rect 14415 5525 14427 5528
rect 14369 5519 14427 5525
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 16853 5559 16911 5565
rect 16853 5525 16865 5559
rect 16899 5556 16911 5559
rect 17144 5556 17172 5596
rect 17494 5584 17500 5596
rect 17552 5584 17558 5636
rect 17954 5624 17960 5636
rect 17915 5596 17960 5624
rect 17954 5584 17960 5596
rect 18012 5584 18018 5636
rect 18230 5584 18236 5636
rect 18288 5624 18294 5636
rect 19334 5624 19340 5636
rect 18288 5596 19340 5624
rect 18288 5584 18294 5596
rect 19334 5584 19340 5596
rect 19392 5624 19398 5636
rect 19705 5627 19763 5633
rect 19705 5624 19717 5627
rect 19392 5596 19717 5624
rect 19392 5584 19398 5596
rect 19705 5593 19717 5596
rect 19751 5593 19763 5627
rect 19705 5587 19763 5593
rect 20254 5584 20260 5636
rect 20312 5624 20318 5636
rect 20533 5627 20591 5633
rect 20533 5624 20545 5627
rect 20312 5596 20545 5624
rect 20312 5584 20318 5596
rect 20533 5593 20545 5596
rect 20579 5593 20591 5627
rect 20533 5587 20591 5593
rect 22278 5584 22284 5636
rect 22336 5624 22342 5636
rect 23658 5624 23664 5636
rect 22336 5596 23664 5624
rect 22336 5584 22342 5596
rect 23658 5584 23664 5596
rect 23716 5584 23722 5636
rect 24857 5627 24915 5633
rect 24857 5593 24869 5627
rect 24903 5624 24915 5627
rect 25038 5624 25044 5636
rect 24903 5596 25044 5624
rect 24903 5593 24915 5596
rect 24857 5587 24915 5593
rect 25038 5584 25044 5596
rect 25096 5624 25102 5636
rect 27338 5624 27344 5636
rect 25096 5596 27344 5624
rect 25096 5584 25102 5596
rect 27338 5584 27344 5596
rect 27396 5584 27402 5636
rect 29178 5584 29184 5636
rect 29236 5624 29242 5636
rect 30662 5627 30720 5633
rect 30662 5624 30674 5627
rect 29236 5596 30674 5624
rect 29236 5584 29242 5596
rect 30662 5593 30674 5596
rect 30708 5593 30720 5627
rect 30760 5624 30788 5664
rect 30929 5661 30941 5695
rect 30975 5692 30987 5695
rect 31478 5692 31484 5704
rect 30975 5664 31484 5692
rect 30975 5661 30987 5664
rect 30929 5655 30987 5661
rect 31478 5652 31484 5664
rect 31536 5652 31542 5704
rect 35894 5652 35900 5704
rect 35952 5692 35958 5704
rect 36173 5695 36231 5701
rect 36173 5692 36185 5695
rect 35952 5664 36185 5692
rect 35952 5652 35958 5664
rect 36173 5661 36185 5664
rect 36219 5661 36231 5695
rect 36173 5655 36231 5661
rect 32582 5624 32588 5636
rect 30760 5596 32588 5624
rect 30662 5587 30720 5593
rect 32582 5584 32588 5596
rect 32640 5624 32646 5636
rect 33045 5627 33103 5633
rect 33045 5624 33057 5627
rect 32640 5596 33057 5624
rect 32640 5584 32646 5596
rect 33045 5593 33057 5596
rect 33091 5593 33103 5627
rect 33045 5587 33103 5593
rect 34790 5584 34796 5636
rect 34848 5624 34854 5636
rect 36970 5627 37028 5633
rect 36970 5624 36982 5627
rect 34848 5596 36982 5624
rect 34848 5584 34854 5596
rect 36970 5593 36982 5596
rect 37016 5593 37028 5627
rect 36970 5587 37028 5593
rect 16899 5528 17172 5556
rect 16899 5525 16911 5528
rect 16853 5519 16911 5525
rect 17218 5516 17224 5568
rect 17276 5556 17282 5568
rect 17773 5559 17831 5565
rect 17773 5556 17785 5559
rect 17276 5528 17785 5556
rect 17276 5516 17282 5528
rect 17773 5525 17785 5528
rect 17819 5525 17831 5559
rect 17773 5519 17831 5525
rect 19426 5516 19432 5568
rect 19484 5556 19490 5568
rect 19797 5559 19855 5565
rect 19797 5556 19809 5559
rect 19484 5528 19809 5556
rect 19484 5516 19490 5528
rect 19797 5525 19809 5528
rect 19843 5525 19855 5559
rect 20714 5556 20720 5568
rect 20675 5528 20720 5556
rect 19797 5519 19855 5525
rect 20714 5516 20720 5528
rect 20772 5516 20778 5568
rect 32490 5556 32496 5568
rect 32451 5528 32496 5556
rect 32490 5516 32496 5528
rect 32548 5516 32554 5568
rect 34514 5516 34520 5568
rect 34572 5556 34578 5568
rect 35069 5559 35127 5565
rect 35069 5556 35081 5559
rect 34572 5528 35081 5556
rect 34572 5516 34578 5528
rect 35069 5525 35081 5528
rect 35115 5525 35127 5559
rect 35069 5519 35127 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 8665 5355 8723 5361
rect 8665 5321 8677 5355
rect 8711 5352 8723 5355
rect 10502 5352 10508 5364
rect 8711 5324 10508 5352
rect 8711 5321 8723 5324
rect 8665 5315 8723 5321
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 10870 5312 10876 5364
rect 10928 5352 10934 5364
rect 10965 5355 11023 5361
rect 10965 5352 10977 5355
rect 10928 5324 10977 5352
rect 10928 5312 10934 5324
rect 10965 5321 10977 5324
rect 11011 5321 11023 5355
rect 15010 5352 15016 5364
rect 10965 5315 11023 5321
rect 13740 5324 15016 5352
rect 10318 5244 10324 5296
rect 10376 5284 10382 5296
rect 13740 5284 13768 5324
rect 15010 5312 15016 5324
rect 15068 5312 15074 5364
rect 15562 5312 15568 5364
rect 15620 5352 15626 5364
rect 15657 5355 15715 5361
rect 15657 5352 15669 5355
rect 15620 5324 15669 5352
rect 15620 5312 15626 5324
rect 15657 5321 15669 5324
rect 15703 5321 15715 5355
rect 19058 5352 19064 5364
rect 19019 5324 19064 5352
rect 15657 5315 15715 5321
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 19978 5312 19984 5364
rect 20036 5352 20042 5364
rect 20349 5355 20407 5361
rect 20349 5352 20361 5355
rect 20036 5324 20361 5352
rect 20036 5312 20042 5324
rect 20349 5321 20361 5324
rect 20395 5352 20407 5355
rect 20714 5352 20720 5364
rect 20395 5324 20720 5352
rect 20395 5321 20407 5324
rect 20349 5315 20407 5321
rect 20714 5312 20720 5324
rect 20772 5312 20778 5364
rect 36633 5355 36691 5361
rect 36633 5352 36645 5355
rect 22066 5324 31754 5352
rect 10376 5256 13768 5284
rect 10376 5244 10382 5256
rect 9674 5176 9680 5228
rect 9732 5216 9738 5228
rect 10597 5219 10655 5225
rect 10597 5216 10609 5219
rect 9732 5188 10609 5216
rect 9732 5176 9738 5188
rect 10597 5185 10609 5188
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 10962 5176 10968 5228
rect 11020 5216 11026 5228
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 11020 5188 11529 5216
rect 11020 5176 11026 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 11698 5216 11704 5228
rect 11659 5188 11704 5216
rect 11517 5179 11575 5185
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 12158 5176 12164 5228
rect 12216 5216 12222 5228
rect 13740 5225 13768 5256
rect 13814 5244 13820 5296
rect 13872 5284 13878 5296
rect 15105 5287 15163 5293
rect 15105 5284 15117 5287
rect 13872 5256 15117 5284
rect 13872 5244 13878 5256
rect 14016 5225 14044 5256
rect 15105 5253 15117 5256
rect 15151 5284 15163 5287
rect 17218 5284 17224 5296
rect 15151 5256 17224 5284
rect 15151 5253 15163 5256
rect 15105 5247 15163 5253
rect 17218 5244 17224 5256
rect 17276 5244 17282 5296
rect 20165 5287 20223 5293
rect 20165 5253 20177 5287
rect 20211 5284 20223 5287
rect 21266 5284 21272 5296
rect 20211 5256 21272 5284
rect 20211 5253 20223 5256
rect 20165 5247 20223 5253
rect 21266 5244 21272 5256
rect 21324 5244 21330 5296
rect 21910 5244 21916 5296
rect 21968 5284 21974 5296
rect 22066 5284 22094 5324
rect 21968 5256 22094 5284
rect 21968 5244 21974 5256
rect 24946 5244 24952 5296
rect 25004 5284 25010 5296
rect 25590 5284 25596 5296
rect 25004 5256 25596 5284
rect 25004 5244 25010 5256
rect 25590 5244 25596 5256
rect 25648 5244 25654 5296
rect 26237 5287 26295 5293
rect 26237 5253 26249 5287
rect 26283 5284 26295 5287
rect 26326 5284 26332 5296
rect 26283 5256 26332 5284
rect 26283 5253 26295 5256
rect 26237 5247 26295 5253
rect 26326 5244 26332 5256
rect 26384 5284 26390 5296
rect 26510 5284 26516 5296
rect 26384 5256 26516 5284
rect 26384 5244 26390 5256
rect 26510 5244 26516 5256
rect 26568 5244 26574 5296
rect 27706 5244 27712 5296
rect 27764 5284 27770 5296
rect 28086 5287 28144 5293
rect 28086 5284 28098 5287
rect 27764 5256 28098 5284
rect 27764 5244 27770 5256
rect 28086 5253 28098 5256
rect 28132 5253 28144 5287
rect 28086 5247 28144 5253
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12216 5188 12909 5216
rect 12216 5176 12222 5188
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 13725 5219 13783 5225
rect 13725 5185 13737 5219
rect 13771 5185 13783 5219
rect 13725 5179 13783 5185
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5185 14059 5219
rect 14001 5179 14059 5185
rect 14185 5219 14243 5225
rect 14185 5185 14197 5219
rect 14231 5216 14243 5219
rect 14829 5219 14887 5225
rect 14829 5216 14841 5219
rect 14231 5188 14841 5216
rect 14231 5185 14243 5188
rect 14185 5179 14243 5185
rect 14829 5185 14841 5188
rect 14875 5216 14887 5219
rect 15562 5216 15568 5228
rect 14875 5188 15056 5216
rect 15523 5188 15568 5216
rect 14875 5185 14887 5188
rect 14829 5179 14887 5185
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10410 5148 10416 5160
rect 10100 5120 10416 5148
rect 10100 5108 10106 5120
rect 10410 5108 10416 5120
rect 10468 5108 10474 5160
rect 12621 5151 12679 5157
rect 12621 5117 12633 5151
rect 12667 5148 12679 5151
rect 12802 5148 12808 5160
rect 12667 5120 12808 5148
rect 12667 5117 12679 5120
rect 12621 5111 12679 5117
rect 12802 5108 12808 5120
rect 12860 5108 12866 5160
rect 13538 5108 13544 5160
rect 13596 5148 13602 5160
rect 13863 5151 13921 5157
rect 13863 5148 13875 5151
rect 13596 5120 13875 5148
rect 13596 5108 13602 5120
rect 13863 5117 13875 5120
rect 13909 5148 13921 5151
rect 14918 5148 14924 5160
rect 13909 5120 14924 5148
rect 13909 5117 13921 5120
rect 13863 5111 13921 5117
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 15028 5148 15056 5188
rect 15562 5176 15568 5188
rect 15620 5176 15626 5228
rect 15654 5176 15660 5228
rect 15712 5216 15718 5228
rect 15841 5219 15899 5225
rect 15841 5216 15853 5219
rect 15712 5188 15853 5216
rect 15712 5176 15718 5188
rect 15841 5185 15853 5188
rect 15887 5216 15899 5219
rect 16390 5216 16396 5228
rect 15887 5188 16396 5216
rect 15887 5185 15899 5188
rect 15841 5179 15899 5185
rect 16390 5176 16396 5188
rect 16448 5176 16454 5228
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5216 16911 5219
rect 16899 5188 17356 5216
rect 16899 5185 16911 5188
rect 16853 5179 16911 5185
rect 16482 5148 16488 5160
rect 15028 5120 16488 5148
rect 16482 5108 16488 5120
rect 16540 5108 16546 5160
rect 17034 5148 17040 5160
rect 16995 5120 17040 5148
rect 17034 5108 17040 5120
rect 17092 5108 17098 5160
rect 17129 5151 17187 5157
rect 17129 5117 17141 5151
rect 17175 5117 17187 5151
rect 17328 5148 17356 5188
rect 17402 5176 17408 5228
rect 17460 5216 17466 5228
rect 18049 5219 18107 5225
rect 18049 5216 18061 5219
rect 17460 5188 18061 5216
rect 17460 5176 17466 5188
rect 18049 5185 18061 5188
rect 18095 5185 18107 5219
rect 18874 5216 18880 5228
rect 18835 5188 18880 5216
rect 18049 5179 18107 5185
rect 18874 5176 18880 5188
rect 18932 5176 18938 5228
rect 19334 5176 19340 5228
rect 19392 5216 19398 5228
rect 19981 5219 20039 5225
rect 19981 5216 19993 5219
rect 19392 5188 19993 5216
rect 19392 5176 19398 5188
rect 19981 5185 19993 5188
rect 20027 5185 20039 5219
rect 19981 5179 20039 5185
rect 20993 5219 21051 5225
rect 20993 5185 21005 5219
rect 21039 5216 21051 5219
rect 24854 5216 24860 5228
rect 21039 5188 24860 5216
rect 21039 5185 21051 5188
rect 20993 5179 21051 5185
rect 24854 5176 24860 5188
rect 24912 5176 24918 5228
rect 25133 5219 25191 5225
rect 25133 5185 25145 5219
rect 25179 5216 25191 5219
rect 27798 5216 27804 5228
rect 25179 5188 27804 5216
rect 25179 5185 25191 5188
rect 25133 5179 25191 5185
rect 27798 5176 27804 5188
rect 27856 5176 27862 5228
rect 17954 5148 17960 5160
rect 17328 5120 17960 5148
rect 17129 5111 17187 5117
rect 7834 5040 7840 5092
rect 7892 5080 7898 5092
rect 9217 5083 9275 5089
rect 9217 5080 9229 5083
rect 7892 5052 9229 5080
rect 7892 5040 7898 5052
rect 9217 5049 9229 5052
rect 9263 5080 9275 5083
rect 10686 5080 10692 5092
rect 9263 5052 10692 5080
rect 9263 5049 9275 5052
rect 9217 5043 9275 5049
rect 10686 5040 10692 5052
rect 10744 5040 10750 5092
rect 12713 5083 12771 5089
rect 12713 5049 12725 5083
rect 12759 5080 12771 5083
rect 16669 5083 16727 5089
rect 16669 5080 16681 5083
rect 12759 5052 16681 5080
rect 12759 5049 12771 5052
rect 12713 5043 12771 5049
rect 16669 5049 16681 5052
rect 16715 5049 16727 5083
rect 17144 5080 17172 5111
rect 17954 5108 17960 5120
rect 18012 5148 18018 5160
rect 23474 5148 23480 5160
rect 18012 5120 22094 5148
rect 23435 5120 23480 5148
rect 18012 5108 18018 5120
rect 17310 5080 17316 5092
rect 17144 5052 17316 5080
rect 16669 5043 16727 5049
rect 17310 5040 17316 5052
rect 17368 5040 17374 5092
rect 18322 5040 18328 5092
rect 18380 5080 18386 5092
rect 20901 5083 20959 5089
rect 20901 5080 20913 5083
rect 18380 5052 20913 5080
rect 18380 5040 18386 5052
rect 20901 5049 20913 5052
rect 20947 5049 20959 5083
rect 22066 5080 22094 5120
rect 23474 5108 23480 5120
rect 23532 5108 23538 5160
rect 28350 5148 28356 5160
rect 28311 5120 28356 5148
rect 28350 5108 28356 5120
rect 28408 5108 28414 5160
rect 31726 5148 31754 5324
rect 32784 5324 36645 5352
rect 32490 5148 32496 5160
rect 31726 5120 32496 5148
rect 32490 5108 32496 5120
rect 32548 5148 32554 5160
rect 32784 5157 32812 5324
rect 36633 5321 36645 5324
rect 36679 5321 36691 5355
rect 36633 5315 36691 5321
rect 32861 5287 32919 5293
rect 32861 5253 32873 5287
rect 32907 5284 32919 5287
rect 33594 5284 33600 5296
rect 32907 5256 33600 5284
rect 32907 5253 32919 5256
rect 32861 5247 32919 5253
rect 33594 5244 33600 5256
rect 33652 5244 33658 5296
rect 33778 5284 33784 5296
rect 33739 5256 33784 5284
rect 33778 5244 33784 5256
rect 33836 5244 33842 5296
rect 35529 5287 35587 5293
rect 35529 5253 35541 5287
rect 35575 5284 35587 5287
rect 36170 5284 36176 5296
rect 35575 5256 36176 5284
rect 35575 5253 35587 5256
rect 35529 5247 35587 5253
rect 36170 5244 36176 5256
rect 36228 5244 36234 5296
rect 36648 5284 36676 5315
rect 36906 5312 36912 5364
rect 36964 5352 36970 5364
rect 37921 5355 37979 5361
rect 37921 5352 37933 5355
rect 36964 5324 37933 5352
rect 36964 5312 36970 5324
rect 37921 5321 37933 5324
rect 37967 5321 37979 5355
rect 37921 5315 37979 5321
rect 37366 5284 37372 5296
rect 36648 5256 37372 5284
rect 37366 5244 37372 5256
rect 37424 5244 37430 5296
rect 35989 5219 36047 5225
rect 35989 5216 36001 5219
rect 33244 5188 36001 5216
rect 32585 5151 32643 5157
rect 32585 5148 32597 5151
rect 32548 5120 32597 5148
rect 32548 5108 32554 5120
rect 32585 5117 32597 5120
rect 32631 5117 32643 5151
rect 32585 5111 32643 5117
rect 32769 5151 32827 5157
rect 32769 5117 32781 5151
rect 32815 5148 32827 5151
rect 32858 5148 32864 5160
rect 32815 5120 32864 5148
rect 32815 5117 32827 5120
rect 32769 5111 32827 5117
rect 26973 5083 27031 5089
rect 26973 5080 26985 5083
rect 22066 5052 26985 5080
rect 20901 5043 20959 5049
rect 26973 5049 26985 5052
rect 27019 5049 27031 5083
rect 29730 5080 29736 5092
rect 26973 5043 27031 5049
rect 28828 5052 29736 5080
rect 7558 5012 7564 5024
rect 7519 4984 7564 5012
rect 7558 4972 7564 4984
rect 7616 4972 7622 5024
rect 8113 5015 8171 5021
rect 8113 4981 8125 5015
rect 8159 5012 8171 5015
rect 9769 5015 9827 5021
rect 9769 5012 9781 5015
rect 8159 4984 9781 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 9769 4981 9781 4984
rect 9815 5012 9827 5015
rect 10502 5012 10508 5024
rect 9815 4984 10508 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 10502 4972 10508 4984
rect 10560 5012 10566 5024
rect 10962 5012 10968 5024
rect 10560 4984 10968 5012
rect 10560 4972 10566 4984
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 11885 5015 11943 5021
rect 11885 4981 11897 5015
rect 11931 5012 11943 5015
rect 12158 5012 12164 5024
rect 11931 4984 12164 5012
rect 11931 4981 11943 4984
rect 11885 4975 11943 4981
rect 12158 4972 12164 4984
rect 12216 4972 12222 5024
rect 13078 5012 13084 5024
rect 13039 4984 13084 5012
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 14093 5015 14151 5021
rect 14093 4981 14105 5015
rect 14139 5012 14151 5015
rect 14182 5012 14188 5024
rect 14139 4984 14188 5012
rect 14139 4981 14151 4984
rect 14093 4975 14151 4981
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 14366 4972 14372 5024
rect 14424 5012 14430 5024
rect 14645 5015 14703 5021
rect 14645 5012 14657 5015
rect 14424 4984 14657 5012
rect 14424 4972 14430 4984
rect 14645 4981 14657 4984
rect 14691 4981 14703 5015
rect 15102 5012 15108 5024
rect 15063 4984 15108 5012
rect 14645 4975 14703 4981
rect 15102 4972 15108 4984
rect 15160 4972 15166 5024
rect 15838 5012 15844 5024
rect 15799 4984 15844 5012
rect 15838 4972 15844 4984
rect 15896 4972 15902 5024
rect 18230 5012 18236 5024
rect 18191 4984 18236 5012
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 21818 5012 21824 5024
rect 21779 4984 21824 5012
rect 21818 4972 21824 4984
rect 21876 4972 21882 5024
rect 28718 4972 28724 5024
rect 28776 5012 28782 5024
rect 28828 5021 28856 5052
rect 29730 5040 29736 5052
rect 29788 5040 29794 5092
rect 32600 5080 32628 5111
rect 32858 5108 32864 5120
rect 32916 5108 32922 5160
rect 33042 5080 33048 5092
rect 32600 5052 33048 5080
rect 33042 5040 33048 5052
rect 33100 5040 33106 5092
rect 33244 5089 33272 5188
rect 35989 5185 36001 5188
rect 36035 5185 36047 5219
rect 37458 5216 37464 5228
rect 37419 5188 37464 5216
rect 35989 5179 36047 5185
rect 37458 5176 37464 5188
rect 37516 5176 37522 5228
rect 38102 5216 38108 5228
rect 38063 5188 38108 5216
rect 38102 5176 38108 5188
rect 38160 5176 38166 5228
rect 33229 5083 33287 5089
rect 33229 5049 33241 5083
rect 33275 5049 33287 5083
rect 33229 5043 33287 5049
rect 36446 5040 36452 5092
rect 36504 5080 36510 5092
rect 37277 5083 37335 5089
rect 37277 5080 37289 5083
rect 36504 5052 37289 5080
rect 36504 5040 36510 5052
rect 37277 5049 37289 5052
rect 37323 5049 37335 5083
rect 37277 5043 37335 5049
rect 28813 5015 28871 5021
rect 28813 5012 28825 5015
rect 28776 4984 28825 5012
rect 28776 4972 28782 4984
rect 28813 4981 28825 4984
rect 28859 4981 28871 5015
rect 29362 5012 29368 5024
rect 29323 4984 29368 5012
rect 28813 4975 28871 4981
rect 29362 4972 29368 4984
rect 29420 4972 29426 5024
rect 29822 4972 29828 5024
rect 29880 5012 29886 5024
rect 29917 5015 29975 5021
rect 29917 5012 29929 5015
rect 29880 4984 29929 5012
rect 29880 4972 29886 4984
rect 29917 4981 29929 4984
rect 29963 4981 29975 5015
rect 30558 5012 30564 5024
rect 30519 4984 30564 5012
rect 29917 4975 29975 4981
rect 30558 4972 30564 4984
rect 30616 4972 30622 5024
rect 31570 5012 31576 5024
rect 31531 4984 31576 5012
rect 31570 4972 31576 4984
rect 31628 4972 31634 5024
rect 36173 5015 36231 5021
rect 36173 4981 36185 5015
rect 36219 5012 36231 5015
rect 36262 5012 36268 5024
rect 36219 4984 36268 5012
rect 36219 4981 36231 4984
rect 36173 4975 36231 4981
rect 36262 4972 36268 4984
rect 36320 4972 36326 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 11701 4811 11759 4817
rect 11701 4777 11713 4811
rect 11747 4808 11759 4811
rect 12618 4808 12624 4820
rect 11747 4780 12624 4808
rect 11747 4777 11759 4780
rect 11701 4771 11759 4777
rect 12618 4768 12624 4780
rect 12676 4808 12682 4820
rect 14461 4811 14519 4817
rect 12676 4780 14412 4808
rect 12676 4768 12682 4780
rect 9398 4740 9404 4752
rect 9311 4712 9404 4740
rect 9398 4700 9404 4712
rect 9456 4740 9462 4752
rect 10597 4743 10655 4749
rect 9456 4712 10272 4740
rect 9456 4700 9462 4712
rect 7837 4675 7895 4681
rect 7837 4641 7849 4675
rect 7883 4672 7895 4675
rect 10134 4672 10140 4684
rect 7883 4644 10140 4672
rect 7883 4641 7895 4644
rect 7837 4635 7895 4641
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 10244 4672 10272 4712
rect 10597 4709 10609 4743
rect 10643 4740 10655 4743
rect 13722 4740 13728 4752
rect 10643 4712 13728 4740
rect 10643 4709 10655 4712
rect 10597 4703 10655 4709
rect 13722 4700 13728 4712
rect 13780 4700 13786 4752
rect 14384 4672 14412 4780
rect 14461 4777 14473 4811
rect 14507 4808 14519 4811
rect 15562 4808 15568 4820
rect 14507 4780 15568 4808
rect 14507 4777 14519 4780
rect 14461 4771 14519 4777
rect 15562 4768 15568 4780
rect 15620 4768 15626 4820
rect 16482 4808 16488 4820
rect 16443 4780 16488 4808
rect 16482 4768 16488 4780
rect 16540 4768 16546 4820
rect 16942 4768 16948 4820
rect 17000 4808 17006 4820
rect 17129 4811 17187 4817
rect 17129 4808 17141 4811
rect 17000 4780 17141 4808
rect 17000 4768 17006 4780
rect 17129 4777 17141 4780
rect 17175 4808 17187 4811
rect 17494 4808 17500 4820
rect 17175 4780 17500 4808
rect 17175 4777 17187 4780
rect 17129 4771 17187 4777
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 17681 4811 17739 4817
rect 17681 4777 17693 4811
rect 17727 4808 17739 4811
rect 19426 4808 19432 4820
rect 17727 4780 19432 4808
rect 17727 4777 17739 4780
rect 17681 4771 17739 4777
rect 19426 4768 19432 4780
rect 19484 4808 19490 4820
rect 20162 4808 20168 4820
rect 19484 4780 20168 4808
rect 19484 4768 19490 4780
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 20254 4768 20260 4820
rect 20312 4808 20318 4820
rect 20349 4811 20407 4817
rect 20349 4808 20361 4811
rect 20312 4780 20361 4808
rect 20312 4768 20318 4780
rect 20349 4777 20361 4780
rect 20395 4777 20407 4811
rect 20349 4771 20407 4777
rect 20993 4811 21051 4817
rect 20993 4777 21005 4811
rect 21039 4808 21051 4811
rect 21082 4808 21088 4820
rect 21039 4780 21088 4808
rect 21039 4777 21051 4780
rect 20993 4771 21051 4777
rect 21082 4768 21088 4780
rect 21140 4768 21146 4820
rect 21266 4768 21272 4820
rect 21324 4808 21330 4820
rect 21324 4780 23704 4808
rect 21324 4768 21330 4780
rect 14918 4700 14924 4752
rect 14976 4740 14982 4752
rect 17034 4740 17040 4752
rect 14976 4712 17040 4740
rect 14976 4700 14982 4712
rect 17034 4700 17040 4712
rect 17092 4700 17098 4752
rect 23676 4740 23704 4780
rect 24578 4768 24584 4820
rect 24636 4808 24642 4820
rect 27065 4811 27123 4817
rect 27065 4808 27077 4811
rect 24636 4780 27077 4808
rect 24636 4768 24642 4780
rect 27065 4777 27077 4780
rect 27111 4777 27123 4811
rect 27065 4771 27123 4777
rect 31849 4811 31907 4817
rect 31849 4777 31861 4811
rect 31895 4808 31907 4811
rect 33686 4808 33692 4820
rect 31895 4780 33692 4808
rect 31895 4777 31907 4780
rect 31849 4771 31907 4777
rect 33686 4768 33692 4780
rect 33744 4768 33750 4820
rect 34149 4811 34207 4817
rect 34149 4777 34161 4811
rect 34195 4808 34207 4811
rect 34514 4808 34520 4820
rect 34195 4780 34520 4808
rect 34195 4777 34207 4780
rect 34149 4771 34207 4777
rect 34514 4768 34520 4780
rect 34572 4768 34578 4820
rect 35437 4811 35495 4817
rect 35437 4777 35449 4811
rect 35483 4808 35495 4811
rect 37458 4808 37464 4820
rect 35483 4780 37464 4808
rect 35483 4777 35495 4780
rect 35437 4771 35495 4777
rect 37458 4768 37464 4780
rect 37516 4768 37522 4820
rect 25225 4743 25283 4749
rect 25225 4740 25237 4743
rect 23676 4712 25237 4740
rect 25225 4709 25237 4712
rect 25271 4709 25283 4743
rect 32030 4740 32036 4752
rect 25225 4703 25283 4709
rect 31220 4712 32036 4740
rect 10244 4644 13124 4672
rect 14384 4644 14504 4672
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4604 7343 4607
rect 9490 4604 9496 4616
rect 7331 4576 9496 4604
rect 7331 4573 7343 4576
rect 7285 4567 7343 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 10410 4604 10416 4616
rect 10371 4576 10416 4604
rect 10410 4564 10416 4576
rect 10468 4564 10474 4616
rect 12710 4604 12716 4616
rect 12671 4576 12716 4604
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 12897 4607 12955 4613
rect 12897 4573 12909 4607
rect 12943 4604 12955 4607
rect 12986 4604 12992 4616
rect 12943 4576 12992 4604
rect 12943 4573 12955 4576
rect 12897 4567 12955 4573
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 13096 4613 13124 4644
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4604 13139 4607
rect 13262 4604 13268 4616
rect 13127 4576 13268 4604
rect 13127 4573 13139 4576
rect 13081 4567 13139 4573
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 14182 4604 14188 4616
rect 14143 4576 14188 4604
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14366 4604 14372 4616
rect 14327 4576 14372 4604
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 14476 4613 14504 4644
rect 15102 4632 15108 4684
rect 15160 4672 15166 4684
rect 18598 4672 18604 4684
rect 15160 4644 18604 4672
rect 15160 4632 15166 4644
rect 18598 4632 18604 4644
rect 18656 4632 18662 4684
rect 31220 4681 31248 4712
rect 32030 4700 32036 4712
rect 32088 4700 32094 4752
rect 35342 4740 35348 4752
rect 34808 4712 35348 4740
rect 30653 4675 30711 4681
rect 22949 4644 24716 4672
rect 14461 4607 14519 4613
rect 14461 4573 14473 4607
rect 14507 4573 14519 4607
rect 14461 4567 14519 4573
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 15654 4604 15660 4616
rect 15427 4576 15660 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 15654 4564 15660 4576
rect 15712 4564 15718 4616
rect 16577 4607 16635 4613
rect 16577 4573 16589 4607
rect 16623 4604 16635 4607
rect 18046 4604 18052 4616
rect 16623 4576 18052 4604
rect 16623 4573 16635 4576
rect 16577 4567 16635 4573
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 18141 4607 18199 4613
rect 18141 4573 18153 4607
rect 18187 4573 18199 4607
rect 18141 4567 18199 4573
rect 6733 4539 6791 4545
rect 6733 4505 6745 4539
rect 6779 4536 6791 4539
rect 8110 4536 8116 4548
rect 6779 4508 8116 4536
rect 6779 4505 6791 4508
rect 6733 4499 6791 4505
rect 8110 4496 8116 4508
rect 8168 4496 8174 4548
rect 8389 4539 8447 4545
rect 8389 4505 8401 4539
rect 8435 4536 8447 4539
rect 11149 4539 11207 4545
rect 8435 4508 11100 4536
rect 8435 4505 8447 4508
rect 8389 4499 8447 4505
rect 5258 4468 5264 4480
rect 5219 4440 5264 4468
rect 5258 4428 5264 4440
rect 5316 4428 5322 4480
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 5905 4471 5963 4477
rect 5905 4468 5917 4471
rect 5684 4440 5917 4468
rect 5684 4428 5690 4440
rect 5905 4437 5917 4440
rect 5951 4437 5963 4471
rect 5905 4431 5963 4437
rect 9953 4471 10011 4477
rect 9953 4437 9965 4471
rect 9999 4468 10011 4471
rect 10962 4468 10968 4480
rect 9999 4440 10968 4468
rect 9999 4437 10011 4440
rect 9953 4431 10011 4437
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 11072 4468 11100 4508
rect 11149 4505 11161 4539
rect 11195 4536 11207 4539
rect 11195 4508 12434 4536
rect 11195 4505 11207 4508
rect 11149 4499 11207 4505
rect 11974 4468 11980 4480
rect 11072 4440 11980 4468
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 12250 4468 12256 4480
rect 12211 4440 12256 4468
rect 12250 4428 12256 4440
rect 12308 4428 12314 4480
rect 12406 4468 12434 4508
rect 15930 4496 15936 4548
rect 15988 4536 15994 4548
rect 18156 4536 18184 4567
rect 19426 4564 19432 4616
rect 19484 4604 19490 4616
rect 19521 4607 19579 4613
rect 19521 4604 19533 4607
rect 19484 4576 19533 4604
rect 19484 4564 19490 4576
rect 19521 4573 19533 4576
rect 19567 4573 19579 4607
rect 19521 4567 19579 4573
rect 20530 4564 20536 4616
rect 20588 4604 20594 4616
rect 22949 4604 22977 4644
rect 20588 4576 22977 4604
rect 23017 4607 23075 4613
rect 20588 4564 20594 4576
rect 23017 4573 23029 4607
rect 23063 4604 23075 4607
rect 23474 4604 23480 4616
rect 23063 4576 23480 4604
rect 23063 4573 23075 4576
rect 23017 4567 23075 4573
rect 23474 4564 23480 4576
rect 23532 4564 23538 4616
rect 23566 4564 23572 4616
rect 23624 4604 23630 4616
rect 24581 4607 24639 4613
rect 24581 4604 24593 4607
rect 23624 4576 24593 4604
rect 23624 4564 23630 4576
rect 24581 4573 24593 4576
rect 24627 4573 24639 4607
rect 24688 4604 24716 4644
rect 30653 4641 30665 4675
rect 30699 4672 30711 4675
rect 31205 4675 31263 4681
rect 31205 4672 31217 4675
rect 30699 4644 31217 4672
rect 30699 4641 30711 4644
rect 30653 4635 30711 4641
rect 31205 4641 31217 4644
rect 31251 4641 31263 4675
rect 31205 4635 31263 4641
rect 31570 4632 31576 4684
rect 31628 4672 31634 4684
rect 31628 4644 32536 4672
rect 31628 4632 31634 4644
rect 26338 4607 26396 4613
rect 26338 4604 26350 4607
rect 24688 4576 26350 4604
rect 24581 4567 24639 4573
rect 26338 4573 26350 4576
rect 26384 4573 26396 4607
rect 26338 4567 26396 4573
rect 26605 4607 26663 4613
rect 26605 4573 26617 4607
rect 26651 4604 26663 4607
rect 27062 4604 27068 4616
rect 26651 4576 27068 4604
rect 26651 4573 26663 4576
rect 26605 4567 26663 4573
rect 27062 4564 27068 4576
rect 27120 4604 27126 4616
rect 28350 4604 28356 4616
rect 27120 4576 28356 4604
rect 27120 4564 27126 4576
rect 28350 4564 28356 4576
rect 28408 4604 28414 4616
rect 28445 4607 28503 4613
rect 28445 4604 28457 4607
rect 28408 4576 28457 4604
rect 28408 4564 28414 4576
rect 28445 4573 28457 4576
rect 28491 4573 28503 4607
rect 28445 4567 28503 4573
rect 30101 4607 30159 4613
rect 30101 4573 30113 4607
rect 30147 4604 30159 4607
rect 32122 4604 32128 4616
rect 30147 4576 32128 4604
rect 30147 4573 30159 4576
rect 30101 4567 30159 4573
rect 32122 4564 32128 4576
rect 32180 4564 32186 4616
rect 32508 4613 32536 4644
rect 33042 4632 33048 4684
rect 33100 4672 33106 4684
rect 34808 4681 34836 4712
rect 35342 4700 35348 4712
rect 35400 4700 35406 4752
rect 37366 4740 37372 4752
rect 37327 4712 37372 4740
rect 37366 4700 37372 4712
rect 37424 4700 37430 4752
rect 34793 4675 34851 4681
rect 34793 4672 34805 4675
rect 33100 4644 34805 4672
rect 33100 4632 33106 4644
rect 34793 4641 34805 4644
rect 34839 4641 34851 4675
rect 34793 4635 34851 4641
rect 34977 4675 35035 4681
rect 34977 4641 34989 4675
rect 35023 4672 35035 4675
rect 35434 4672 35440 4684
rect 35023 4644 35440 4672
rect 35023 4641 35035 4644
rect 34977 4635 35035 4641
rect 35434 4632 35440 4644
rect 35492 4632 35498 4684
rect 32493 4607 32551 4613
rect 32493 4573 32505 4607
rect 32539 4573 32551 4607
rect 32493 4567 32551 4573
rect 32674 4564 32680 4616
rect 32732 4604 32738 4616
rect 32950 4604 32956 4616
rect 32732 4576 32956 4604
rect 32732 4564 32738 4576
rect 32950 4564 32956 4576
rect 33008 4564 33014 4616
rect 33870 4564 33876 4616
rect 33928 4604 33934 4616
rect 33965 4607 34023 4613
rect 33965 4604 33977 4607
rect 33928 4576 33977 4604
rect 33928 4564 33934 4576
rect 33965 4573 33977 4576
rect 34011 4604 34023 4607
rect 34054 4604 34060 4616
rect 34011 4576 34060 4604
rect 34011 4573 34023 4576
rect 33965 4567 34023 4573
rect 34054 4564 34060 4576
rect 34112 4564 34118 4616
rect 35989 4607 36047 4613
rect 35989 4573 36001 4607
rect 36035 4604 36047 4607
rect 36078 4604 36084 4616
rect 36035 4576 36084 4604
rect 36035 4573 36047 4576
rect 35989 4567 36047 4573
rect 36078 4564 36084 4576
rect 36136 4564 36142 4616
rect 36262 4613 36268 4616
rect 36256 4604 36268 4613
rect 36223 4576 36268 4604
rect 36256 4567 36268 4576
rect 36262 4564 36268 4567
rect 36320 4564 36326 4616
rect 37918 4564 37924 4616
rect 37976 4604 37982 4616
rect 38105 4607 38163 4613
rect 38105 4604 38117 4607
rect 37976 4576 38117 4604
rect 37976 4564 37982 4576
rect 38105 4573 38117 4576
rect 38151 4573 38163 4607
rect 38105 4567 38163 4573
rect 15988 4508 18184 4536
rect 19720 4508 21772 4536
rect 15988 4496 15994 4508
rect 15194 4468 15200 4480
rect 12406 4440 15200 4468
rect 15194 4428 15200 4440
rect 15252 4428 15258 4480
rect 15841 4471 15899 4477
rect 15841 4437 15853 4471
rect 15887 4468 15899 4471
rect 16850 4468 16856 4480
rect 15887 4440 16856 4468
rect 15887 4437 15899 4440
rect 15841 4431 15899 4437
rect 16850 4428 16856 4440
rect 16908 4428 16914 4480
rect 18325 4471 18383 4477
rect 18325 4437 18337 4471
rect 18371 4468 18383 4471
rect 19242 4468 19248 4480
rect 18371 4440 19248 4468
rect 18371 4437 18383 4440
rect 18325 4431 18383 4437
rect 19242 4428 19248 4440
rect 19300 4428 19306 4480
rect 19720 4477 19748 4508
rect 19705 4471 19763 4477
rect 19705 4437 19717 4471
rect 19751 4437 19763 4471
rect 19705 4431 19763 4437
rect 20438 4428 20444 4480
rect 20496 4468 20502 4480
rect 21266 4468 21272 4480
rect 20496 4440 21272 4468
rect 20496 4428 20502 4440
rect 21266 4428 21272 4440
rect 21324 4428 21330 4480
rect 21634 4468 21640 4480
rect 21595 4440 21640 4468
rect 21634 4428 21640 4440
rect 21692 4428 21698 4480
rect 21744 4468 21772 4508
rect 22370 4496 22376 4548
rect 22428 4536 22434 4548
rect 22750 4539 22808 4545
rect 22750 4536 22762 4539
rect 22428 4508 22762 4536
rect 22428 4496 22434 4508
rect 22750 4505 22762 4508
rect 22796 4505 22808 4539
rect 22750 4499 22808 4505
rect 23661 4539 23719 4545
rect 23661 4505 23673 4539
rect 23707 4536 23719 4539
rect 23842 4536 23848 4548
rect 23707 4508 23848 4536
rect 23707 4505 23719 4508
rect 23661 4499 23719 4505
rect 23842 4496 23848 4508
rect 23900 4496 23906 4548
rect 26418 4496 26424 4548
rect 26476 4536 26482 4548
rect 28178 4539 28236 4545
rect 28178 4536 28190 4539
rect 26476 4508 28190 4536
rect 26476 4496 26482 4508
rect 28178 4505 28190 4508
rect 28224 4505 28236 4539
rect 28178 4499 28236 4505
rect 31202 4496 31208 4548
rect 31260 4536 31266 4548
rect 31389 4539 31447 4545
rect 31389 4536 31401 4539
rect 31260 4508 31401 4536
rect 31260 4496 31266 4508
rect 31389 4505 31401 4508
rect 31435 4505 31447 4539
rect 31389 4499 31447 4505
rect 31481 4539 31539 4545
rect 31481 4505 31493 4539
rect 31527 4536 31539 4539
rect 31527 4508 32352 4536
rect 31527 4505 31539 4508
rect 31481 4499 31539 4505
rect 22094 4468 22100 4480
rect 21744 4440 22100 4468
rect 22094 4428 22100 4440
rect 22152 4428 22158 4480
rect 24765 4471 24823 4477
rect 24765 4437 24777 4471
rect 24811 4468 24823 4471
rect 27154 4468 27160 4480
rect 24811 4440 27160 4468
rect 24811 4437 24823 4440
rect 24765 4431 24823 4437
rect 27154 4428 27160 4440
rect 27212 4428 27218 4480
rect 28994 4468 29000 4480
rect 28955 4440 29000 4468
rect 28994 4428 29000 4440
rect 29052 4428 29058 4480
rect 29914 4468 29920 4480
rect 29875 4440 29920 4468
rect 29914 4428 29920 4440
rect 29972 4428 29978 4480
rect 32324 4477 32352 4508
rect 36538 4496 36544 4548
rect 36596 4536 36602 4548
rect 36596 4508 37964 4536
rect 36596 4496 36602 4508
rect 32309 4471 32367 4477
rect 32309 4437 32321 4471
rect 32355 4437 32367 4471
rect 33134 4468 33140 4480
rect 33095 4440 33140 4468
rect 32309 4431 32367 4437
rect 33134 4428 33140 4440
rect 33192 4428 33198 4480
rect 35066 4428 35072 4480
rect 35124 4468 35130 4480
rect 37936 4477 37964 4508
rect 37921 4471 37979 4477
rect 35124 4440 35169 4468
rect 35124 4428 35130 4440
rect 37921 4437 37933 4471
rect 37967 4437 37979 4471
rect 37921 4431 37979 4437
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 8297 4267 8355 4273
rect 8297 4233 8309 4267
rect 8343 4264 8355 4267
rect 8570 4264 8576 4276
rect 8343 4236 8576 4264
rect 8343 4233 8355 4236
rect 8297 4227 8355 4233
rect 8570 4224 8576 4236
rect 8628 4264 8634 4276
rect 9398 4264 9404 4276
rect 8628 4236 9404 4264
rect 8628 4224 8634 4236
rect 9398 4224 9404 4236
rect 9456 4224 9462 4276
rect 10410 4224 10416 4276
rect 10468 4264 10474 4276
rect 10597 4267 10655 4273
rect 10597 4264 10609 4267
rect 10468 4236 10609 4264
rect 10468 4224 10474 4236
rect 10597 4233 10609 4236
rect 10643 4233 10655 4267
rect 10597 4227 10655 4233
rect 10686 4224 10692 4276
rect 10744 4264 10750 4276
rect 12986 4264 12992 4276
rect 10744 4236 12992 4264
rect 10744 4224 10750 4236
rect 12986 4224 12992 4236
rect 13044 4224 13050 4276
rect 15654 4224 15660 4276
rect 15712 4264 15718 4276
rect 17770 4264 17776 4276
rect 15712 4236 17776 4264
rect 15712 4224 15718 4236
rect 17770 4224 17776 4236
rect 17828 4224 17834 4276
rect 18414 4224 18420 4276
rect 18472 4264 18478 4276
rect 23566 4264 23572 4276
rect 18472 4236 23572 4264
rect 18472 4224 18478 4236
rect 23566 4224 23572 4236
rect 23624 4224 23630 4276
rect 28442 4264 28448 4276
rect 28403 4236 28448 4264
rect 28442 4224 28448 4236
rect 28500 4224 28506 4276
rect 28905 4267 28963 4273
rect 28905 4233 28917 4267
rect 28951 4233 28963 4267
rect 28905 4227 28963 4233
rect 12894 4196 12900 4208
rect 10060 4168 10364 4196
rect 7745 4131 7803 4137
rect 7745 4097 7757 4131
rect 7791 4128 7803 4131
rect 10060 4128 10088 4168
rect 10226 4128 10232 4140
rect 7791 4100 10088 4128
rect 10187 4100 10232 4128
rect 7791 4097 7803 4100
rect 7745 4091 7803 4097
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 10336 4128 10364 4168
rect 12544 4168 12900 4196
rect 11514 4128 11520 4140
rect 10336 4100 11520 4128
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 12066 4128 12072 4140
rect 12027 4100 12072 4128
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12434 4088 12440 4140
rect 12492 4128 12498 4140
rect 12544 4128 12572 4168
rect 12894 4156 12900 4168
rect 12952 4156 12958 4208
rect 13280 4168 14136 4196
rect 12710 4128 12716 4140
rect 12492 4100 12572 4128
rect 12671 4100 12716 4128
rect 12492 4088 12498 4100
rect 12710 4088 12716 4100
rect 12768 4088 12774 4140
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 9030 4060 9036 4072
rect 6687 4032 9036 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 10042 4060 10048 4072
rect 10003 4032 10048 4060
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 10137 4063 10195 4069
rect 10137 4029 10149 4063
rect 10183 4060 10195 4063
rect 10410 4060 10416 4072
rect 10183 4032 10416 4060
rect 10183 4029 10195 4032
rect 10137 4023 10195 4029
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 11609 4063 11667 4069
rect 11609 4029 11621 4063
rect 11655 4060 11667 4063
rect 13280 4060 13308 4168
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4097 13415 4131
rect 13538 4128 13544 4140
rect 13499 4100 13544 4128
rect 13357 4091 13415 4097
rect 11655 4032 13308 4060
rect 13372 4060 13400 4091
rect 13538 4088 13544 4100
rect 13596 4088 13602 4140
rect 13722 4088 13728 4140
rect 13780 4128 13786 4140
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13780 4100 14013 4128
rect 13780 4088 13786 4100
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 13814 4060 13820 4072
rect 13372 4032 13820 4060
rect 11655 4029 11667 4032
rect 11609 4023 11667 4029
rect 13814 4020 13820 4032
rect 13872 4020 13878 4072
rect 14108 4060 14136 4168
rect 16482 4156 16488 4208
rect 16540 4196 16546 4208
rect 19705 4199 19763 4205
rect 19705 4196 19717 4199
rect 16540 4168 19717 4196
rect 16540 4156 16546 4168
rect 19705 4165 19717 4168
rect 19751 4165 19763 4199
rect 21082 4196 21088 4208
rect 19705 4159 19763 4165
rect 19904 4168 21088 4196
rect 14734 4088 14740 4140
rect 14792 4128 14798 4140
rect 15562 4128 15568 4140
rect 14792 4100 15568 4128
rect 14792 4088 14798 4100
rect 15562 4088 15568 4100
rect 15620 4128 15626 4140
rect 15657 4131 15715 4137
rect 15657 4128 15669 4131
rect 15620 4100 15669 4128
rect 15620 4088 15626 4100
rect 15657 4097 15669 4100
rect 15703 4097 15715 4131
rect 16850 4128 16856 4140
rect 15657 4091 15715 4097
rect 15764 4100 16856 4128
rect 15764 4060 15792 4100
rect 16850 4088 16856 4100
rect 16908 4088 16914 4140
rect 17218 4128 17224 4140
rect 17179 4100 17224 4128
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 17586 4128 17592 4140
rect 17547 4100 17592 4128
rect 17586 4088 17592 4100
rect 17644 4088 17650 4140
rect 17770 4128 17776 4140
rect 17731 4100 17776 4128
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 18049 4131 18107 4137
rect 18049 4097 18061 4131
rect 18095 4097 18107 4131
rect 18049 4091 18107 4097
rect 18233 4131 18291 4137
rect 18233 4097 18245 4131
rect 18279 4128 18291 4131
rect 18322 4128 18328 4140
rect 18279 4100 18328 4128
rect 18279 4097 18291 4100
rect 18233 4091 18291 4097
rect 14108 4032 15792 4060
rect 15838 4020 15844 4072
rect 15896 4060 15902 4072
rect 16390 4060 16396 4072
rect 15896 4032 16396 4060
rect 15896 4020 15902 4032
rect 16390 4020 16396 4032
rect 16448 4060 16454 4072
rect 17954 4060 17960 4072
rect 16448 4032 17960 4060
rect 16448 4020 16454 4032
rect 17954 4020 17960 4032
rect 18012 4020 18018 4072
rect 5813 3995 5871 4001
rect 5813 3961 5825 3995
rect 5859 3992 5871 3995
rect 7282 3992 7288 4004
rect 5859 3964 7288 3992
rect 5859 3961 5871 3964
rect 5813 3955 5871 3961
rect 7282 3952 7288 3964
rect 7340 3952 7346 4004
rect 8849 3995 8907 4001
rect 8849 3961 8861 3995
rect 8895 3992 8907 3995
rect 10594 3992 10600 4004
rect 8895 3964 10600 3992
rect 8895 3961 8907 3964
rect 8849 3955 8907 3961
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 12434 3992 12440 4004
rect 10704 3964 12440 3992
rect 3973 3927 4031 3933
rect 3973 3893 3985 3927
rect 4019 3924 4031 3927
rect 4062 3924 4068 3936
rect 4019 3896 4068 3924
rect 4019 3893 4031 3896
rect 3973 3887 4031 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4614 3924 4620 3936
rect 4575 3896 4620 3924
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 5261 3927 5319 3933
rect 5261 3893 5273 3927
rect 5307 3924 5319 3927
rect 5534 3924 5540 3936
rect 5307 3896 5540 3924
rect 5307 3893 5319 3896
rect 5261 3887 5319 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 7190 3924 7196 3936
rect 7151 3896 7196 3924
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 9398 3924 9404 3936
rect 9359 3896 9404 3924
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 9582 3884 9588 3936
rect 9640 3924 9646 3936
rect 10704 3924 10732 3964
rect 12434 3952 12440 3964
rect 12492 3952 12498 4004
rect 12802 3952 12808 4004
rect 12860 3992 12866 4004
rect 13357 3995 13415 4001
rect 13357 3992 13369 3995
rect 12860 3964 13369 3992
rect 12860 3952 12866 3964
rect 13357 3961 13369 3964
rect 13403 3961 13415 3995
rect 14274 3992 14280 4004
rect 13357 3955 13415 3961
rect 13832 3964 14280 3992
rect 12250 3924 12256 3936
rect 9640 3896 10732 3924
rect 12211 3896 12256 3924
rect 9640 3884 9646 3896
rect 12250 3884 12256 3896
rect 12308 3884 12314 3936
rect 12897 3927 12955 3933
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 13832 3924 13860 3964
rect 14274 3952 14280 3964
rect 14332 3952 14338 4004
rect 15197 3995 15255 4001
rect 15197 3961 15209 3995
rect 15243 3992 15255 3995
rect 15746 3992 15752 4004
rect 15243 3964 15752 3992
rect 15243 3961 15255 3964
rect 15197 3955 15255 3961
rect 15746 3952 15752 3964
rect 15804 3952 15810 4004
rect 18064 3992 18092 4091
rect 18322 4088 18328 4100
rect 18380 4088 18386 4140
rect 18693 4131 18751 4137
rect 18693 4097 18705 4131
rect 18739 4128 18751 4131
rect 19334 4128 19340 4140
rect 18739 4100 19340 4128
rect 18739 4097 18751 4100
rect 18693 4091 18751 4097
rect 19334 4088 19340 4100
rect 19392 4128 19398 4140
rect 19613 4131 19671 4137
rect 19392 4100 19472 4128
rect 19392 4088 19398 4100
rect 19444 4069 19472 4100
rect 19613 4097 19625 4131
rect 19659 4128 19671 4131
rect 19904 4128 19932 4168
rect 21082 4156 21088 4168
rect 21140 4156 21146 4208
rect 23934 4156 23940 4208
rect 23992 4196 23998 4208
rect 28920 4196 28948 4227
rect 31202 4224 31208 4276
rect 31260 4264 31266 4276
rect 31481 4267 31539 4273
rect 31481 4264 31493 4267
rect 31260 4236 31493 4264
rect 31260 4224 31266 4236
rect 31481 4233 31493 4236
rect 31527 4264 31539 4267
rect 31662 4264 31668 4276
rect 31527 4236 31668 4264
rect 31527 4233 31539 4236
rect 31481 4227 31539 4233
rect 31662 4224 31668 4236
rect 31720 4224 31726 4276
rect 32122 4264 32128 4276
rect 32083 4236 32128 4264
rect 32122 4224 32128 4236
rect 32180 4224 32186 4276
rect 33134 4224 33140 4276
rect 33192 4264 33198 4276
rect 33781 4267 33839 4273
rect 33781 4264 33793 4267
rect 33192 4236 33793 4264
rect 33192 4224 33198 4236
rect 33781 4233 33793 4236
rect 33827 4233 33839 4267
rect 33781 4227 33839 4233
rect 34793 4267 34851 4273
rect 34793 4233 34805 4267
rect 34839 4264 34851 4267
rect 35066 4264 35072 4276
rect 34839 4236 35072 4264
rect 34839 4233 34851 4236
rect 34793 4227 34851 4233
rect 35066 4224 35072 4236
rect 35124 4224 35130 4276
rect 35345 4267 35403 4273
rect 35345 4233 35357 4267
rect 35391 4264 35403 4267
rect 35434 4264 35440 4276
rect 35391 4236 35440 4264
rect 35391 4233 35403 4236
rect 35345 4227 35403 4233
rect 35434 4224 35440 4236
rect 35492 4224 35498 4276
rect 23992 4168 28948 4196
rect 29816 4199 29874 4205
rect 23992 4156 23998 4168
rect 29816 4165 29828 4199
rect 29862 4196 29874 4199
rect 29914 4196 29920 4208
rect 29862 4168 29920 4196
rect 29862 4165 29874 4168
rect 29816 4159 29874 4165
rect 29914 4156 29920 4168
rect 29972 4156 29978 4208
rect 32490 4196 32496 4208
rect 32451 4168 32496 4196
rect 32490 4156 32496 4168
rect 32548 4156 32554 4208
rect 33042 4156 33048 4208
rect 33100 4196 33106 4208
rect 33100 4168 33180 4196
rect 33100 4156 33106 4168
rect 19659 4100 19932 4128
rect 19659 4097 19671 4100
rect 19613 4091 19671 4097
rect 19978 4088 19984 4140
rect 20036 4128 20042 4140
rect 20533 4131 20591 4137
rect 20533 4128 20545 4131
rect 20036 4100 20545 4128
rect 20036 4088 20042 4100
rect 20533 4097 20545 4100
rect 20579 4097 20591 4131
rect 21174 4128 21180 4140
rect 21135 4100 21180 4128
rect 20533 4091 20591 4097
rect 21174 4088 21180 4100
rect 21232 4088 21238 4140
rect 21266 4088 21272 4140
rect 21324 4128 21330 4140
rect 22738 4128 22744 4140
rect 21324 4100 22744 4128
rect 21324 4088 21330 4100
rect 22738 4088 22744 4100
rect 22796 4128 22802 4140
rect 22925 4131 22983 4137
rect 22925 4128 22937 4131
rect 22796 4100 22937 4128
rect 22796 4088 22802 4100
rect 22925 4097 22937 4100
rect 22971 4097 22983 4131
rect 22925 4091 22983 4097
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 24121 4131 24179 4137
rect 24121 4128 24133 4131
rect 23532 4100 24133 4128
rect 23532 4088 23538 4100
rect 24121 4097 24133 4100
rect 24167 4097 24179 4131
rect 24121 4091 24179 4097
rect 24210 4088 24216 4140
rect 24268 4128 24274 4140
rect 24377 4131 24435 4137
rect 24377 4128 24389 4131
rect 24268 4100 24389 4128
rect 24268 4088 24274 4100
rect 24377 4097 24389 4100
rect 24423 4097 24435 4131
rect 24377 4091 24435 4097
rect 27154 4088 27160 4140
rect 27212 4128 27218 4140
rect 27321 4131 27379 4137
rect 27321 4128 27333 4131
rect 27212 4100 27333 4128
rect 27212 4088 27218 4100
rect 27321 4097 27333 4100
rect 27367 4097 27379 4131
rect 27321 4091 27379 4097
rect 28258 4088 28264 4140
rect 28316 4128 28322 4140
rect 28994 4128 29000 4140
rect 28316 4100 29000 4128
rect 28316 4088 28322 4100
rect 28994 4088 29000 4100
rect 29052 4128 29058 4140
rect 29089 4131 29147 4137
rect 29089 4128 29101 4131
rect 29052 4100 29101 4128
rect 29052 4088 29058 4100
rect 29089 4097 29101 4100
rect 29135 4097 29147 4131
rect 32582 4128 32588 4140
rect 29089 4091 29147 4097
rect 31726 4100 32588 4128
rect 19429 4063 19487 4069
rect 19429 4029 19441 4063
rect 19475 4029 19487 4063
rect 24026 4060 24032 4072
rect 19429 4023 19487 4029
rect 19720 4032 24032 4060
rect 19720 3992 19748 4032
rect 24026 4020 24032 4032
rect 24084 4020 24090 4072
rect 27062 4060 27068 4072
rect 27023 4032 27068 4060
rect 27062 4020 27068 4032
rect 27120 4020 27126 4072
rect 28442 4020 28448 4072
rect 28500 4060 28506 4072
rect 29549 4063 29607 4069
rect 29549 4060 29561 4063
rect 28500 4032 29561 4060
rect 28500 4020 28506 4032
rect 29549 4029 29561 4032
rect 29595 4029 29607 4063
rect 29549 4023 29607 4029
rect 20070 3992 20076 4004
rect 18064 3964 19748 3992
rect 20031 3964 20076 3992
rect 20070 3952 20076 3964
rect 20128 3952 20134 4004
rect 20162 3952 20168 4004
rect 20220 3992 20226 4004
rect 21818 3992 21824 4004
rect 20220 3964 21824 3992
rect 20220 3952 20226 3964
rect 21818 3952 21824 3964
rect 21876 3952 21882 4004
rect 26053 3995 26111 4001
rect 22066 3964 23244 3992
rect 12943 3896 13860 3924
rect 14185 3927 14243 3933
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 14185 3893 14197 3927
rect 14231 3924 14243 3927
rect 14366 3924 14372 3936
rect 14231 3896 14372 3924
rect 14231 3893 14243 3896
rect 14185 3887 14243 3893
rect 14366 3884 14372 3896
rect 14424 3924 14430 3936
rect 15470 3924 15476 3936
rect 14424 3896 15476 3924
rect 14424 3884 14430 3896
rect 15470 3884 15476 3896
rect 15528 3884 15534 3936
rect 15838 3924 15844 3936
rect 15799 3896 15844 3924
rect 15838 3884 15844 3896
rect 15896 3884 15902 3936
rect 16758 3924 16764 3936
rect 16719 3896 16764 3924
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 20717 3927 20775 3933
rect 20717 3893 20729 3927
rect 20763 3924 20775 3927
rect 21082 3924 21088 3936
rect 20763 3896 21088 3924
rect 20763 3893 20775 3896
rect 20717 3887 20775 3893
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 21266 3884 21272 3936
rect 21324 3924 21330 3936
rect 22066 3924 22094 3964
rect 23216 3936 23244 3964
rect 26053 3961 26065 3995
rect 26099 3992 26111 3995
rect 26234 3992 26240 4004
rect 26099 3964 26240 3992
rect 26099 3961 26111 3964
rect 26053 3955 26111 3961
rect 26234 3952 26240 3964
rect 26292 3992 26298 4004
rect 26970 3992 26976 4004
rect 26292 3964 26976 3992
rect 26292 3952 26298 3964
rect 26970 3952 26976 3964
rect 27028 3952 27034 4004
rect 30929 3995 30987 4001
rect 30929 3961 30941 3995
rect 30975 3992 30987 3995
rect 31726 3992 31754 4100
rect 32582 4088 32588 4100
rect 32640 4088 32646 4140
rect 32030 4020 32036 4072
rect 32088 4060 32094 4072
rect 32677 4063 32735 4069
rect 32677 4060 32689 4063
rect 32088 4032 32689 4060
rect 32088 4020 32094 4032
rect 32677 4029 32689 4032
rect 32723 4060 32735 4063
rect 33042 4060 33048 4072
rect 32723 4032 33048 4060
rect 32723 4029 32735 4032
rect 32677 4023 32735 4029
rect 33042 4020 33048 4032
rect 33100 4020 33106 4072
rect 33152 4060 33180 4168
rect 36078 4156 36084 4208
rect 36136 4196 36142 4208
rect 36354 4196 36360 4208
rect 36136 4168 36360 4196
rect 36136 4156 36142 4168
rect 36354 4156 36360 4168
rect 36412 4196 36418 4208
rect 36412 4168 36768 4196
rect 36412 4156 36418 4168
rect 33226 4088 33232 4140
rect 33284 4128 33290 4140
rect 34609 4131 34667 4137
rect 34609 4128 34621 4131
rect 33284 4100 34621 4128
rect 33284 4088 33290 4100
rect 34609 4097 34621 4100
rect 34655 4128 34667 4131
rect 35986 4128 35992 4140
rect 34655 4100 35992 4128
rect 34655 4097 34667 4100
rect 34609 4091 34667 4097
rect 35986 4088 35992 4100
rect 36044 4088 36050 4140
rect 36446 4088 36452 4140
rect 36504 4137 36510 4140
rect 36740 4137 36768 4168
rect 36504 4128 36516 4137
rect 36725 4131 36783 4137
rect 36504 4100 36549 4128
rect 36504 4091 36516 4100
rect 36725 4097 36737 4131
rect 36771 4097 36783 4131
rect 37461 4131 37519 4137
rect 37461 4128 37473 4131
rect 36725 4091 36783 4097
rect 36832 4100 37473 4128
rect 36504 4088 36510 4091
rect 33505 4063 33563 4069
rect 33505 4060 33517 4063
rect 33152 4032 33517 4060
rect 33505 4029 33517 4032
rect 33551 4029 33563 4063
rect 33505 4023 33563 4029
rect 33689 4063 33747 4069
rect 33689 4029 33701 4063
rect 33735 4060 33747 4063
rect 35710 4060 35716 4072
rect 33735 4032 35716 4060
rect 33735 4029 33747 4032
rect 33689 4023 33747 4029
rect 35710 4020 35716 4032
rect 35768 4020 35774 4072
rect 30975 3964 31754 3992
rect 34149 3995 34207 4001
rect 30975 3961 30987 3964
rect 30929 3955 30987 3961
rect 34149 3961 34161 3995
rect 34195 3992 34207 3995
rect 34195 3964 35848 3992
rect 34195 3961 34207 3964
rect 34149 3955 34207 3961
rect 22462 3924 22468 3936
rect 21324 3896 22094 3924
rect 22375 3896 22468 3924
rect 21324 3884 21330 3896
rect 22462 3884 22468 3896
rect 22520 3924 22526 3936
rect 22830 3924 22836 3936
rect 22520 3896 22836 3924
rect 22520 3884 22526 3896
rect 22830 3884 22836 3896
rect 22888 3884 22894 3936
rect 23198 3884 23204 3936
rect 23256 3924 23262 3936
rect 23477 3927 23535 3933
rect 23477 3924 23489 3927
rect 23256 3896 23489 3924
rect 23256 3884 23262 3896
rect 23477 3893 23489 3896
rect 23523 3893 23535 3927
rect 25498 3924 25504 3936
rect 25459 3896 25504 3924
rect 23477 3887 23535 3893
rect 25498 3884 25504 3896
rect 25556 3884 25562 3936
rect 28534 3884 28540 3936
rect 28592 3924 28598 3936
rect 29454 3924 29460 3936
rect 28592 3896 29460 3924
rect 28592 3884 28598 3896
rect 29454 3884 29460 3896
rect 29512 3884 29518 3936
rect 35820 3924 35848 3964
rect 36832 3924 36860 4100
rect 37461 4097 37473 4100
rect 37507 4097 37519 4131
rect 37461 4091 37519 4097
rect 37734 4088 37740 4140
rect 37792 4128 37798 4140
rect 38105 4131 38163 4137
rect 38105 4128 38117 4131
rect 37792 4100 38117 4128
rect 37792 4088 37798 4100
rect 38105 4097 38117 4100
rect 38151 4097 38163 4131
rect 38105 4091 38163 4097
rect 37182 3952 37188 4004
rect 37240 3992 37246 4004
rect 37921 3995 37979 4001
rect 37921 3992 37933 3995
rect 37240 3964 37933 3992
rect 37240 3952 37246 3964
rect 37921 3961 37933 3964
rect 37967 3961 37979 3995
rect 37921 3955 37979 3961
rect 37274 3924 37280 3936
rect 35820 3896 36860 3924
rect 37235 3896 37280 3924
rect 37274 3884 37280 3896
rect 37332 3884 37338 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 7834 3720 7840 3732
rect 7524 3692 7840 3720
rect 7524 3680 7530 3692
rect 7834 3680 7840 3692
rect 7892 3680 7898 3732
rect 8389 3723 8447 3729
rect 8389 3689 8401 3723
rect 8435 3720 8447 3723
rect 8754 3720 8760 3732
rect 8435 3692 8760 3720
rect 8435 3689 8447 3692
rect 8389 3683 8447 3689
rect 8754 3680 8760 3692
rect 8812 3720 8818 3732
rect 9582 3720 9588 3732
rect 8812 3692 9588 3720
rect 8812 3680 8818 3692
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 10226 3680 10232 3732
rect 10284 3720 10290 3732
rect 10321 3723 10379 3729
rect 10321 3720 10333 3723
rect 10284 3692 10333 3720
rect 10284 3680 10290 3692
rect 10321 3689 10333 3692
rect 10367 3689 10379 3723
rect 10321 3683 10379 3689
rect 11701 3723 11759 3729
rect 11701 3689 11713 3723
rect 11747 3720 11759 3723
rect 13446 3720 13452 3732
rect 11747 3692 13452 3720
rect 11747 3689 11759 3692
rect 11701 3683 11759 3689
rect 13446 3680 13452 3692
rect 13504 3680 13510 3732
rect 14366 3720 14372 3732
rect 14327 3692 14372 3720
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 16574 3680 16580 3732
rect 16632 3720 16638 3732
rect 16669 3723 16727 3729
rect 16669 3720 16681 3723
rect 16632 3692 16681 3720
rect 16632 3680 16638 3692
rect 16669 3689 16681 3692
rect 16715 3720 16727 3723
rect 17126 3720 17132 3732
rect 16715 3692 17132 3720
rect 16715 3689 16727 3692
rect 16669 3683 16727 3689
rect 17126 3680 17132 3692
rect 17184 3680 17190 3732
rect 18325 3723 18383 3729
rect 18325 3689 18337 3723
rect 18371 3720 18383 3723
rect 18414 3720 18420 3732
rect 18371 3692 18420 3720
rect 18371 3689 18383 3692
rect 18325 3683 18383 3689
rect 18414 3680 18420 3692
rect 18472 3680 18478 3732
rect 18874 3680 18880 3732
rect 18932 3720 18938 3732
rect 19245 3723 19303 3729
rect 19245 3720 19257 3723
rect 18932 3692 19257 3720
rect 18932 3680 18938 3692
rect 19245 3689 19257 3692
rect 19291 3689 19303 3723
rect 19245 3683 19303 3689
rect 19334 3680 19340 3732
rect 19392 3720 19398 3732
rect 22738 3720 22744 3732
rect 19392 3692 22600 3720
rect 22699 3692 22744 3720
rect 19392 3680 19398 3692
rect 6178 3652 6184 3664
rect 6139 3624 6184 3652
rect 6178 3612 6184 3624
rect 6236 3612 6242 3664
rect 7285 3655 7343 3661
rect 7285 3621 7297 3655
rect 7331 3652 7343 3655
rect 12618 3652 12624 3664
rect 7331 3624 12624 3652
rect 7331 3621 7343 3624
rect 7285 3615 7343 3621
rect 12618 3612 12624 3624
rect 12676 3612 12682 3664
rect 13262 3652 13268 3664
rect 12728 3624 13268 3652
rect 6733 3587 6791 3593
rect 6733 3553 6745 3587
rect 6779 3584 6791 3587
rect 11698 3584 11704 3596
rect 6779 3556 11704 3584
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 4062 3516 4068 3528
rect 4023 3488 4068 3516
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3516 5687 3519
rect 8202 3516 8208 3528
rect 5675 3488 8208 3516
rect 5675 3485 5687 3488
rect 5629 3479 5687 3485
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3516 9183 3519
rect 9582 3516 9588 3528
rect 9171 3488 9588 3516
rect 9171 3485 9183 3488
rect 9125 3479 9183 3485
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10134 3516 10140 3528
rect 10095 3488 10140 3516
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 10888 3525 10916 3556
rect 11698 3544 11704 3556
rect 11756 3544 11762 3596
rect 12158 3584 12164 3596
rect 12119 3556 12164 3584
rect 12158 3544 12164 3556
rect 12216 3544 12222 3596
rect 12728 3584 12756 3624
rect 13262 3612 13268 3624
rect 13320 3612 13326 3664
rect 14645 3655 14703 3661
rect 14645 3621 14657 3655
rect 14691 3652 14703 3655
rect 15289 3655 15347 3661
rect 15289 3652 15301 3655
rect 14691 3624 15301 3652
rect 14691 3621 14703 3624
rect 14645 3615 14703 3621
rect 15289 3621 15301 3624
rect 15335 3621 15347 3655
rect 15289 3615 15347 3621
rect 15381 3655 15439 3661
rect 15381 3621 15393 3655
rect 15427 3652 15439 3655
rect 15654 3652 15660 3664
rect 15427 3624 15660 3652
rect 15427 3621 15439 3624
rect 15381 3615 15439 3621
rect 15654 3612 15660 3624
rect 15712 3612 15718 3664
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 21266 3652 21272 3664
rect 20772 3624 21272 3652
rect 20772 3612 20778 3624
rect 21266 3612 21272 3624
rect 21324 3612 21330 3664
rect 22572 3652 22600 3692
rect 22738 3680 22744 3692
rect 22796 3680 22802 3732
rect 23014 3680 23020 3732
rect 23072 3720 23078 3732
rect 26418 3720 26424 3732
rect 23072 3692 26424 3720
rect 23072 3680 23078 3692
rect 26418 3680 26424 3692
rect 26476 3680 26482 3732
rect 26513 3723 26571 3729
rect 26513 3689 26525 3723
rect 26559 3720 26571 3723
rect 27062 3720 27068 3732
rect 26559 3692 27068 3720
rect 26559 3689 26571 3692
rect 26513 3683 26571 3689
rect 27062 3680 27068 3692
rect 27120 3680 27126 3732
rect 28994 3720 29000 3732
rect 28955 3692 29000 3720
rect 28994 3680 29000 3692
rect 29052 3680 29058 3732
rect 29086 3680 29092 3732
rect 29144 3720 29150 3732
rect 30098 3720 30104 3732
rect 29144 3692 30104 3720
rect 29144 3680 29150 3692
rect 30098 3680 30104 3692
rect 30156 3680 30162 3732
rect 33594 3680 33600 3732
rect 33652 3720 33658 3732
rect 36817 3723 36875 3729
rect 36817 3720 36829 3723
rect 33652 3692 36829 3720
rect 33652 3680 33658 3692
rect 36817 3689 36829 3692
rect 36863 3689 36875 3723
rect 36817 3683 36875 3689
rect 28261 3655 28319 3661
rect 28261 3652 28273 3655
rect 22572 3624 28273 3652
rect 28261 3621 28273 3624
rect 28307 3621 28319 3655
rect 28261 3615 28319 3621
rect 28442 3612 28448 3664
rect 28500 3652 28506 3664
rect 34977 3655 35035 3661
rect 34977 3652 34989 3655
rect 28500 3624 34989 3652
rect 28500 3612 28506 3624
rect 34977 3621 34989 3624
rect 35023 3621 35035 3655
rect 34977 3615 35035 3621
rect 36538 3612 36544 3664
rect 36596 3652 36602 3664
rect 38102 3652 38108 3664
rect 36596 3624 38108 3652
rect 36596 3612 36602 3624
rect 38102 3612 38108 3624
rect 38160 3612 38166 3664
rect 12406 3556 12756 3584
rect 10873 3519 10931 3525
rect 10873 3485 10885 3519
rect 10919 3485 10931 3519
rect 11146 3516 11152 3528
rect 10873 3479 10931 3485
rect 10980 3488 11152 3516
rect 5077 3451 5135 3457
rect 5077 3417 5089 3451
rect 5123 3448 5135 3451
rect 6822 3448 6828 3460
rect 5123 3420 6828 3448
rect 5123 3417 5135 3420
rect 5077 3411 5135 3417
rect 6822 3408 6828 3420
rect 6880 3408 6886 3460
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 10980 3448 11008 3488
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 11514 3516 11520 3528
rect 11475 3488 11520 3516
rect 11514 3476 11520 3488
rect 11572 3476 11578 3528
rect 12406 3525 12434 3556
rect 12986 3544 12992 3596
rect 13044 3584 13050 3596
rect 14369 3587 14427 3593
rect 13044 3556 13584 3584
rect 13044 3544 13050 3556
rect 12406 3519 12470 3525
rect 12406 3488 12424 3519
rect 12412 3485 12424 3488
rect 12458 3485 12470 3519
rect 12529 3519 12587 3525
rect 12529 3506 12541 3519
rect 12575 3506 12587 3519
rect 12621 3519 12679 3525
rect 12412 3479 12470 3485
rect 6972 3420 11008 3448
rect 11072 3420 11836 3448
rect 6972 3408 6978 3420
rect 2866 3340 2872 3392
rect 2924 3380 2930 3392
rect 3145 3383 3203 3389
rect 3145 3380 3157 3383
rect 2924 3352 3157 3380
rect 2924 3340 2930 3352
rect 3145 3349 3157 3352
rect 3191 3349 3203 3383
rect 3145 3343 3203 3349
rect 4249 3383 4307 3389
rect 4249 3349 4261 3383
rect 4295 3380 4307 3383
rect 4890 3380 4896 3392
rect 4295 3352 4896 3380
rect 4295 3349 4307 3352
rect 4249 3343 4307 3349
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 9306 3380 9312 3392
rect 9267 3352 9312 3380
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 10870 3380 10876 3392
rect 10100 3352 10876 3380
rect 10100 3340 10106 3352
rect 10870 3340 10876 3352
rect 10928 3340 10934 3392
rect 11072 3389 11100 3420
rect 11057 3383 11115 3389
rect 11057 3349 11069 3383
rect 11103 3349 11115 3383
rect 11808 3380 11836 3420
rect 11882 3408 11888 3460
rect 11940 3448 11946 3460
rect 12299 3451 12357 3457
rect 12526 3454 12532 3506
rect 12584 3454 12590 3506
rect 12621 3485 12633 3519
rect 12667 3516 12679 3519
rect 12667 3488 12848 3516
rect 12667 3485 12679 3488
rect 12621 3479 12679 3485
rect 12299 3448 12311 3451
rect 11940 3420 12311 3448
rect 11940 3408 11946 3420
rect 12299 3417 12311 3420
rect 12345 3417 12357 3451
rect 12820 3448 12848 3488
rect 12894 3476 12900 3528
rect 12952 3516 12958 3528
rect 13556 3525 13584 3556
rect 14369 3553 14381 3587
rect 14415 3584 14427 3587
rect 14550 3584 14556 3596
rect 14415 3556 14556 3584
rect 14415 3553 14427 3556
rect 14369 3547 14427 3553
rect 14550 3544 14556 3556
rect 14608 3544 14614 3596
rect 14826 3544 14832 3596
rect 14884 3584 14890 3596
rect 16482 3584 16488 3596
rect 14884 3556 16488 3584
rect 14884 3544 14890 3556
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 16850 3544 16856 3596
rect 16908 3584 16914 3596
rect 17681 3587 17739 3593
rect 17681 3584 17693 3587
rect 16908 3556 17693 3584
rect 16908 3544 16914 3556
rect 17681 3553 17693 3556
rect 17727 3553 17739 3587
rect 19702 3584 19708 3596
rect 19663 3556 19708 3584
rect 17681 3547 17739 3553
rect 19702 3544 19708 3556
rect 19760 3544 19766 3596
rect 19889 3587 19947 3593
rect 19889 3553 19901 3587
rect 19935 3584 19947 3587
rect 20162 3584 20168 3596
rect 19935 3556 20168 3584
rect 19935 3553 19947 3556
rect 19889 3547 19947 3553
rect 20162 3544 20168 3556
rect 20220 3544 20226 3596
rect 21082 3544 21088 3596
rect 21140 3584 21146 3596
rect 26234 3584 26240 3596
rect 21140 3556 21496 3584
rect 21140 3544 21146 3556
rect 13357 3519 13415 3525
rect 13357 3516 13369 3519
rect 12952 3488 13369 3516
rect 12952 3476 12958 3488
rect 13357 3485 13369 3488
rect 13403 3485 13415 3519
rect 13357 3479 13415 3485
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3485 13599 3519
rect 14458 3516 14464 3528
rect 14419 3488 14464 3516
rect 13541 3479 13599 3485
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3485 15439 3519
rect 16390 3516 16396 3528
rect 16351 3488 16396 3516
rect 15381 3479 15439 3485
rect 13449 3451 13507 3457
rect 13449 3448 13461 3451
rect 12820 3420 13461 3448
rect 12299 3411 12357 3417
rect 13449 3417 13461 3420
rect 13495 3417 13507 3451
rect 13449 3411 13507 3417
rect 14185 3451 14243 3457
rect 14185 3417 14197 3451
rect 14231 3448 14243 3451
rect 14274 3448 14280 3460
rect 14231 3420 14280 3448
rect 14231 3417 14243 3420
rect 14185 3411 14243 3417
rect 14274 3408 14280 3420
rect 14332 3408 14338 3460
rect 15102 3448 15108 3460
rect 15063 3420 15108 3448
rect 15102 3408 15108 3420
rect 15160 3408 15166 3460
rect 12526 3380 12532 3392
rect 11808 3352 12532 3380
rect 11057 3343 11115 3349
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 12805 3383 12863 3389
rect 12805 3349 12817 3383
rect 12851 3380 12863 3383
rect 13722 3380 13728 3392
rect 12851 3352 13728 3380
rect 12851 3349 12863 3352
rect 12805 3343 12863 3349
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 13814 3340 13820 3392
rect 13872 3380 13878 3392
rect 15286 3380 15292 3392
rect 13872 3352 15292 3380
rect 13872 3340 13878 3352
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 15396 3380 15424 3479
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 17865 3519 17923 3525
rect 17865 3516 17877 3519
rect 16816 3488 17877 3516
rect 16816 3476 16822 3488
rect 17865 3485 17877 3488
rect 17911 3516 17923 3519
rect 20530 3516 20536 3528
rect 17911 3488 20536 3516
rect 17911 3485 17923 3488
rect 17865 3479 17923 3485
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 20717 3519 20775 3525
rect 20717 3485 20729 3519
rect 20763 3516 20775 3519
rect 21174 3516 21180 3528
rect 20763 3488 21180 3516
rect 20763 3485 20775 3488
rect 20717 3479 20775 3485
rect 21174 3476 21180 3488
rect 21232 3476 21238 3528
rect 21358 3516 21364 3528
rect 21319 3488 21364 3516
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 21468 3516 21496 3556
rect 24688 3556 26240 3584
rect 21617 3519 21675 3525
rect 21617 3516 21629 3519
rect 21468 3488 21629 3516
rect 21617 3485 21629 3488
rect 21663 3485 21675 3519
rect 21617 3479 21675 3485
rect 23477 3519 23535 3525
rect 23477 3485 23489 3519
rect 23523 3516 23535 3519
rect 23842 3516 23848 3528
rect 23523 3488 23848 3516
rect 23523 3485 23535 3488
rect 23477 3479 23535 3485
rect 23842 3476 23848 3488
rect 23900 3516 23906 3528
rect 24578 3516 24584 3528
rect 23900 3488 24584 3516
rect 23900 3476 23906 3488
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 24688 3525 24716 3556
rect 26234 3544 26240 3556
rect 26292 3544 26298 3596
rect 26418 3544 26424 3596
rect 26476 3584 26482 3596
rect 26878 3584 26884 3596
rect 26476 3556 26884 3584
rect 26476 3544 26482 3556
rect 26878 3544 26884 3556
rect 26936 3544 26942 3596
rect 27154 3544 27160 3596
rect 27212 3584 27218 3596
rect 27212 3556 28488 3584
rect 27212 3544 27218 3556
rect 24673 3519 24731 3525
rect 24673 3485 24685 3519
rect 24719 3485 24731 3519
rect 24673 3479 24731 3485
rect 24762 3476 24768 3528
rect 24820 3516 24826 3528
rect 25409 3519 25467 3525
rect 24820 3488 25360 3516
rect 24820 3476 24826 3488
rect 16666 3448 16672 3460
rect 16627 3420 16672 3448
rect 16666 3408 16672 3420
rect 16724 3408 16730 3460
rect 17957 3451 18015 3457
rect 17957 3417 17969 3451
rect 18003 3448 18015 3451
rect 23934 3448 23940 3460
rect 18003 3420 23940 3448
rect 18003 3417 18015 3420
rect 17957 3411 18015 3417
rect 23934 3408 23940 3420
rect 23992 3408 23998 3460
rect 16209 3383 16267 3389
rect 16209 3380 16221 3383
rect 15396 3352 16221 3380
rect 16209 3349 16221 3352
rect 16255 3349 16267 3383
rect 16209 3343 16267 3349
rect 16298 3340 16304 3392
rect 16356 3380 16362 3392
rect 19613 3383 19671 3389
rect 19613 3380 19625 3383
rect 16356 3352 19625 3380
rect 16356 3340 16362 3352
rect 19613 3349 19625 3352
rect 19659 3349 19671 3383
rect 19613 3343 19671 3349
rect 20070 3340 20076 3392
rect 20128 3380 20134 3392
rect 20533 3383 20591 3389
rect 20533 3380 20545 3383
rect 20128 3352 20545 3380
rect 20128 3340 20134 3352
rect 20533 3349 20545 3352
rect 20579 3349 20591 3383
rect 20533 3343 20591 3349
rect 22830 3340 22836 3392
rect 22888 3380 22894 3392
rect 23293 3383 23351 3389
rect 23293 3380 23305 3383
rect 22888 3352 23305 3380
rect 22888 3340 22894 3352
rect 23293 3349 23305 3352
rect 23339 3349 23351 3383
rect 23293 3343 23351 3349
rect 23842 3340 23848 3392
rect 23900 3380 23906 3392
rect 24489 3383 24547 3389
rect 24489 3380 24501 3383
rect 23900 3352 24501 3380
rect 23900 3340 23906 3352
rect 24489 3349 24501 3352
rect 24535 3349 24547 3383
rect 24489 3343 24547 3349
rect 24946 3340 24952 3392
rect 25004 3380 25010 3392
rect 25225 3383 25283 3389
rect 25225 3380 25237 3383
rect 25004 3352 25237 3380
rect 25004 3340 25010 3352
rect 25225 3349 25237 3352
rect 25271 3349 25283 3383
rect 25332 3380 25360 3488
rect 25409 3485 25421 3519
rect 25455 3516 25467 3519
rect 25590 3516 25596 3528
rect 25455 3488 25596 3516
rect 25455 3485 25467 3488
rect 25409 3479 25467 3485
rect 25590 3476 25596 3488
rect 25648 3476 25654 3528
rect 27798 3516 27804 3528
rect 27759 3488 27804 3516
rect 27798 3476 27804 3488
rect 27856 3476 27862 3528
rect 28460 3525 28488 3556
rect 33042 3544 33048 3596
rect 33100 3584 33106 3596
rect 33505 3587 33563 3593
rect 33505 3584 33517 3587
rect 33100 3556 33517 3584
rect 33100 3544 33106 3556
rect 33505 3553 33517 3556
rect 33551 3553 33563 3587
rect 36354 3584 36360 3596
rect 36315 3556 36360 3584
rect 33505 3547 33563 3553
rect 36354 3544 36360 3556
rect 36412 3544 36418 3596
rect 37734 3584 37740 3596
rect 36464 3556 37740 3584
rect 28445 3519 28503 3525
rect 28445 3485 28457 3519
rect 28491 3516 28503 3519
rect 29549 3519 29607 3525
rect 29549 3516 29561 3519
rect 28491 3488 29561 3516
rect 28491 3485 28503 3488
rect 28445 3479 28503 3485
rect 29549 3485 29561 3488
rect 29595 3485 29607 3519
rect 32953 3519 33011 3525
rect 32953 3516 32965 3519
rect 29549 3479 29607 3485
rect 31726 3488 32965 3516
rect 27816 3448 27844 3476
rect 31726 3448 31754 3488
rect 32953 3485 32965 3488
rect 32999 3516 33011 3519
rect 33778 3516 33784 3528
rect 32999 3488 33784 3516
rect 32999 3485 33011 3488
rect 32953 3479 33011 3485
rect 33778 3476 33784 3488
rect 33836 3476 33842 3528
rect 35342 3476 35348 3528
rect 35400 3516 35406 3528
rect 36464 3516 36492 3556
rect 37734 3544 37740 3556
rect 37792 3544 37798 3596
rect 36998 3516 37004 3528
rect 35400 3488 36492 3516
rect 36959 3488 37004 3516
rect 35400 3476 35406 3488
rect 36998 3476 37004 3488
rect 37056 3476 37062 3528
rect 37642 3516 37648 3528
rect 37603 3488 37648 3516
rect 37642 3476 37648 3488
rect 37700 3476 37706 3528
rect 27816 3420 31754 3448
rect 32214 3408 32220 3460
rect 32272 3448 32278 3460
rect 35986 3448 35992 3460
rect 32272 3420 35992 3448
rect 32272 3408 32278 3420
rect 35986 3408 35992 3420
rect 36044 3408 36050 3460
rect 36112 3451 36170 3457
rect 36112 3417 36124 3451
rect 36158 3448 36170 3451
rect 37550 3448 37556 3460
rect 36158 3420 37556 3448
rect 36158 3417 36170 3420
rect 36112 3411 36170 3417
rect 37550 3408 37556 3420
rect 37608 3408 37614 3460
rect 28442 3380 28448 3392
rect 25332 3352 28448 3380
rect 25225 3343 25283 3349
rect 28442 3340 28448 3352
rect 28500 3340 28506 3392
rect 30190 3340 30196 3392
rect 30248 3380 30254 3392
rect 30653 3383 30711 3389
rect 30653 3380 30665 3383
rect 30248 3352 30665 3380
rect 30248 3340 30254 3352
rect 30653 3349 30665 3352
rect 30699 3349 30711 3383
rect 31478 3380 31484 3392
rect 31439 3352 31484 3380
rect 30653 3343 30711 3349
rect 31478 3340 31484 3352
rect 31536 3340 31542 3392
rect 33410 3340 33416 3392
rect 33468 3380 33474 3392
rect 33594 3380 33600 3392
rect 33468 3352 33600 3380
rect 33468 3340 33474 3352
rect 33594 3340 33600 3352
rect 33652 3380 33658 3392
rect 33689 3383 33747 3389
rect 33689 3380 33701 3383
rect 33652 3352 33701 3380
rect 33652 3340 33658 3352
rect 33689 3349 33701 3352
rect 33735 3349 33747 3383
rect 33689 3343 33747 3349
rect 33778 3340 33784 3392
rect 33836 3380 33842 3392
rect 34149 3383 34207 3389
rect 33836 3352 33881 3380
rect 33836 3340 33842 3352
rect 34149 3349 34161 3383
rect 34195 3380 34207 3383
rect 34790 3380 34796 3392
rect 34195 3352 34796 3380
rect 34195 3349 34207 3352
rect 34149 3343 34207 3349
rect 34790 3340 34796 3352
rect 34848 3340 34854 3392
rect 35802 3340 35808 3392
rect 35860 3380 35866 3392
rect 37461 3383 37519 3389
rect 37461 3380 37473 3383
rect 35860 3352 37473 3380
rect 35860 3340 35866 3352
rect 37461 3349 37473 3352
rect 37507 3349 37519 3383
rect 37461 3343 37519 3349
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 5810 3176 5816 3188
rect 5771 3148 5816 3176
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 7006 3176 7012 3188
rect 6967 3148 7012 3176
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 7745 3179 7803 3185
rect 7745 3145 7757 3179
rect 7791 3176 7803 3179
rect 9217 3179 9275 3185
rect 9217 3176 9229 3179
rect 7791 3148 9229 3176
rect 7791 3145 7803 3148
rect 7745 3139 7803 3145
rect 9217 3145 9229 3148
rect 9263 3145 9275 3179
rect 9582 3176 9588 3188
rect 9543 3148 9588 3176
rect 9217 3139 9275 3145
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 12526 3136 12532 3188
rect 12584 3176 12590 3188
rect 13630 3176 13636 3188
rect 12584 3148 13636 3176
rect 12584 3136 12590 3148
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 14001 3179 14059 3185
rect 14001 3145 14013 3179
rect 14047 3176 14059 3179
rect 15102 3176 15108 3188
rect 14047 3148 15108 3176
rect 14047 3145 14059 3148
rect 14001 3139 14059 3145
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 15565 3179 15623 3185
rect 15565 3145 15577 3179
rect 15611 3176 15623 3179
rect 15930 3176 15936 3188
rect 15611 3148 15792 3176
rect 15891 3148 15936 3176
rect 15611 3145 15623 3148
rect 15565 3139 15623 3145
rect 3053 3111 3111 3117
rect 3053 3077 3065 3111
rect 3099 3108 3111 3111
rect 6914 3108 6920 3120
rect 3099 3080 6920 3108
rect 3099 3077 3111 3080
rect 3053 3071 3111 3077
rect 3804 3049 3832 3080
rect 6914 3068 6920 3080
rect 6972 3068 6978 3120
rect 9030 3068 9036 3120
rect 9088 3108 9094 3120
rect 11882 3108 11888 3120
rect 9088 3080 10548 3108
rect 9088 3068 9094 3080
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3009 3847 3043
rect 3789 3003 3847 3009
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 4614 3040 4620 3052
rect 4387 3012 4620 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3040 5043 3043
rect 5074 3040 5080 3052
rect 5031 3012 5080 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5074 3000 5080 3012
rect 5132 3040 5138 3052
rect 5258 3040 5264 3052
rect 5132 3012 5264 3040
rect 5132 3000 5138 3012
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 5626 3040 5632 3052
rect 5587 3012 5632 3040
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 6822 3040 6828 3052
rect 6783 3012 6828 3040
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 7558 3040 7564 3052
rect 7519 3012 7564 3040
rect 7558 3000 7564 3012
rect 7616 3040 7622 3052
rect 7834 3040 7840 3052
rect 7616 3012 7840 3040
rect 7616 3000 7622 3012
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 8110 3000 8116 3052
rect 8168 3040 8174 3052
rect 8205 3043 8263 3049
rect 8205 3040 8217 3043
rect 8168 3012 8217 3040
rect 8168 3000 8174 3012
rect 8205 3009 8217 3012
rect 8251 3040 8263 3043
rect 8846 3040 8852 3052
rect 8251 3012 8852 3040
rect 8251 3009 8263 3012
rect 8205 3003 8263 3009
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 10042 3040 10048 3052
rect 9048 3012 10048 3040
rect 9048 2981 9076 3012
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 10226 3040 10232 3052
rect 10187 3012 10232 3040
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 10520 3040 10548 3080
rect 10796 3080 11888 3108
rect 10686 3040 10692 3052
rect 10520 3012 10692 3040
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 9033 2975 9091 2981
rect 9033 2941 9045 2975
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 9122 2932 9128 2984
rect 9180 2972 9186 2984
rect 10321 2975 10379 2981
rect 9180 2944 9225 2972
rect 9180 2932 9186 2944
rect 10321 2941 10333 2975
rect 10367 2941 10379 2975
rect 10321 2935 10379 2941
rect 10597 2975 10655 2981
rect 10597 2941 10609 2975
rect 10643 2972 10655 2975
rect 10796 2972 10824 3080
rect 11882 3068 11888 3080
rect 11940 3068 11946 3120
rect 15764 3108 15792 3148
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 17402 3176 17408 3188
rect 17363 3148 17408 3176
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 17586 3136 17592 3188
rect 17644 3176 17650 3188
rect 17865 3179 17923 3185
rect 17865 3176 17877 3179
rect 17644 3148 17877 3176
rect 17644 3136 17650 3148
rect 17865 3145 17877 3148
rect 17911 3145 17923 3179
rect 19978 3176 19984 3188
rect 19939 3148 19984 3176
rect 17865 3139 17923 3145
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 23014 3176 23020 3188
rect 20272 3148 23020 3176
rect 19334 3108 19340 3120
rect 15764 3080 19340 3108
rect 19334 3068 19340 3080
rect 19392 3068 19398 3120
rect 20162 3108 20168 3120
rect 19444 3080 20168 3108
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 11848 3012 11989 3040
rect 11848 3000 11854 3012
rect 11977 3009 11989 3012
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 12989 3044 13047 3049
rect 12989 3043 13124 3044
rect 12989 3009 13001 3043
rect 13035 3016 13124 3043
rect 13035 3009 13047 3016
rect 12989 3003 13047 3009
rect 10643 2944 10824 2972
rect 10643 2941 10655 2944
rect 10597 2935 10655 2941
rect 4525 2907 4583 2913
rect 4525 2873 4537 2907
rect 4571 2904 4583 2907
rect 9950 2904 9956 2916
rect 4571 2876 9956 2904
rect 4571 2873 4583 2876
rect 4525 2867 4583 2873
rect 9950 2864 9956 2876
rect 10008 2864 10014 2916
rect 10336 2904 10364 2935
rect 10870 2932 10876 2984
rect 10928 2972 10934 2984
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 10928 2944 11713 2972
rect 10928 2932 10934 2944
rect 11701 2941 11713 2944
rect 11747 2941 11759 2975
rect 11882 2972 11888 2984
rect 11843 2944 11888 2972
rect 11701 2935 11759 2941
rect 11882 2932 11888 2944
rect 11940 2932 11946 2984
rect 12802 2972 12808 2984
rect 11992 2944 12808 2972
rect 11992 2904 12020 2944
rect 12802 2932 12808 2944
rect 12860 2932 12866 2984
rect 10336 2876 12020 2904
rect 1762 2836 1768 2848
rect 1723 2808 1768 2836
rect 1762 2796 1768 2808
rect 1820 2796 1826 2848
rect 2314 2836 2320 2848
rect 2275 2808 2320 2836
rect 2314 2796 2320 2808
rect 2372 2796 2378 2848
rect 3418 2796 3424 2848
rect 3476 2836 3482 2848
rect 3605 2839 3663 2845
rect 3605 2836 3617 2839
rect 3476 2808 3617 2836
rect 3476 2796 3482 2808
rect 3605 2805 3617 2808
rect 3651 2805 3663 2839
rect 5166 2836 5172 2848
rect 5127 2808 5172 2836
rect 3605 2799 3663 2805
rect 5166 2796 5172 2808
rect 5224 2796 5230 2848
rect 8386 2836 8392 2848
rect 8347 2808 8392 2836
rect 8386 2796 8392 2808
rect 8444 2796 8450 2848
rect 12345 2839 12403 2845
rect 12345 2805 12357 2839
rect 12391 2836 12403 2839
rect 13096 2836 13124 3016
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3040 13691 3043
rect 13814 3040 13820 3052
rect 13679 3012 13820 3040
rect 13679 3009 13691 3012
rect 13633 3003 13691 3009
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 13998 3000 14004 3052
rect 14056 3040 14062 3052
rect 14553 3043 14611 3049
rect 14553 3040 14565 3043
rect 14056 3012 14565 3040
rect 14056 3000 14062 3012
rect 14553 3009 14565 3012
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 15304 3012 15608 3040
rect 13446 2932 13452 2984
rect 13504 2972 13510 2984
rect 13725 2975 13783 2981
rect 13725 2972 13737 2975
rect 13504 2944 13737 2972
rect 13504 2932 13510 2944
rect 13725 2941 13737 2944
rect 13771 2941 13783 2975
rect 14568 2972 14596 3003
rect 15304 2981 15332 3012
rect 15289 2975 15347 2981
rect 14568 2944 15240 2972
rect 13725 2935 13783 2941
rect 13173 2907 13231 2913
rect 13173 2873 13185 2907
rect 13219 2904 13231 2907
rect 15102 2904 15108 2916
rect 13219 2876 15108 2904
rect 13219 2873 13231 2876
rect 13173 2867 13231 2873
rect 15102 2864 15108 2876
rect 15160 2864 15166 2916
rect 13630 2836 13636 2848
rect 12391 2808 13124 2836
rect 13591 2808 13636 2836
rect 12391 2805 12403 2808
rect 12345 2799 12403 2805
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 14734 2836 14740 2848
rect 14695 2808 14740 2836
rect 14734 2796 14740 2808
rect 14792 2796 14798 2848
rect 15212 2836 15240 2944
rect 15289 2941 15301 2975
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 15378 2932 15384 2984
rect 15436 2972 15442 2984
rect 15473 2975 15531 2981
rect 15473 2972 15485 2975
rect 15436 2944 15485 2972
rect 15436 2932 15442 2944
rect 15473 2941 15485 2944
rect 15519 2941 15531 2975
rect 15580 2972 15608 3012
rect 15746 3000 15752 3052
rect 15804 3040 15810 3052
rect 16942 3040 16948 3052
rect 15804 3012 16948 3040
rect 15804 3000 15810 3012
rect 16942 3000 16948 3012
rect 17000 3000 17006 3052
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 17862 3040 17868 3052
rect 17083 3012 17868 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 17862 3000 17868 3012
rect 17920 3000 17926 3052
rect 18138 3040 18144 3052
rect 18099 3012 18144 3040
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 16850 2972 16856 2984
rect 15580 2944 16856 2972
rect 15473 2935 15531 2941
rect 15488 2904 15516 2935
rect 16850 2932 16856 2944
rect 16908 2932 16914 2984
rect 17494 2932 17500 2984
rect 17552 2972 17558 2984
rect 18432 2972 18460 3003
rect 18782 2972 18788 2984
rect 17552 2944 18788 2972
rect 17552 2932 17558 2944
rect 18782 2932 18788 2944
rect 18840 2932 18846 2984
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 19444 2981 19472 3080
rect 20162 3068 20168 3080
rect 20220 3068 20226 3120
rect 19610 3040 19616 3052
rect 19571 3012 19616 3040
rect 19610 3000 19616 3012
rect 19668 3000 19674 3052
rect 19429 2975 19487 2981
rect 19429 2972 19441 2975
rect 19392 2944 19441 2972
rect 19392 2932 19398 2944
rect 19429 2941 19441 2944
rect 19475 2941 19487 2975
rect 19429 2935 19487 2941
rect 19521 2975 19579 2981
rect 19521 2941 19533 2975
rect 19567 2972 19579 2975
rect 20162 2972 20168 2984
rect 19567 2944 20168 2972
rect 19567 2941 19579 2944
rect 19521 2935 19579 2941
rect 20162 2932 20168 2944
rect 20220 2932 20226 2984
rect 20272 2904 20300 3148
rect 23014 3136 23020 3148
rect 23072 3136 23078 3188
rect 23198 3176 23204 3188
rect 23159 3148 23204 3176
rect 23198 3136 23204 3148
rect 23256 3136 23262 3188
rect 24026 3136 24032 3188
rect 24084 3176 24090 3188
rect 25866 3176 25872 3188
rect 24084 3148 25452 3176
rect 25827 3148 25872 3176
rect 24084 3136 24090 3148
rect 23474 3108 23480 3120
rect 21836 3080 23480 3108
rect 20901 3043 20959 3049
rect 20901 3009 20913 3043
rect 20947 3040 20959 3043
rect 20990 3040 20996 3052
rect 20947 3012 20996 3040
rect 20947 3009 20959 3012
rect 20901 3003 20959 3009
rect 20990 3000 20996 3012
rect 21048 3000 21054 3052
rect 21358 3000 21364 3052
rect 21416 3040 21422 3052
rect 21836 3049 21864 3080
rect 23474 3068 23480 3080
rect 23532 3108 23538 3120
rect 24118 3108 24124 3120
rect 23532 3080 24124 3108
rect 23532 3068 23538 3080
rect 24118 3068 24124 3080
rect 24176 3068 24182 3120
rect 25424 3108 25452 3148
rect 25866 3136 25872 3148
rect 25924 3136 25930 3188
rect 28813 3179 28871 3185
rect 28813 3176 28825 3179
rect 25976 3148 28825 3176
rect 25976 3108 26004 3148
rect 28813 3145 28825 3148
rect 28859 3145 28871 3179
rect 30834 3176 30840 3188
rect 30795 3148 30840 3176
rect 28813 3139 28871 3145
rect 30834 3136 30840 3148
rect 30892 3136 30898 3188
rect 31573 3179 31631 3185
rect 31573 3145 31585 3179
rect 31619 3176 31631 3179
rect 33778 3176 33784 3188
rect 31619 3148 33784 3176
rect 31619 3145 31631 3148
rect 31573 3139 31631 3145
rect 33778 3136 33784 3148
rect 33836 3136 33842 3188
rect 33962 3176 33968 3188
rect 33923 3148 33968 3176
rect 33962 3136 33968 3148
rect 34020 3136 34026 3188
rect 35069 3179 35127 3185
rect 35069 3145 35081 3179
rect 35115 3176 35127 3179
rect 35710 3176 35716 3188
rect 35115 3148 35716 3176
rect 35115 3145 35127 3148
rect 35069 3139 35127 3145
rect 35710 3136 35716 3148
rect 35768 3136 35774 3188
rect 35986 3136 35992 3188
rect 36044 3176 36050 3188
rect 37918 3176 37924 3188
rect 36044 3148 37924 3176
rect 36044 3136 36050 3148
rect 37918 3136 37924 3148
rect 37976 3136 37982 3188
rect 25424 3080 26004 3108
rect 26421 3111 26479 3117
rect 26421 3077 26433 3111
rect 26467 3108 26479 3111
rect 27430 3108 27436 3120
rect 26467 3080 27436 3108
rect 26467 3077 26479 3080
rect 26421 3071 26479 3077
rect 22094 3049 22100 3052
rect 21821 3043 21879 3049
rect 21821 3040 21833 3043
rect 21416 3012 21833 3040
rect 21416 3000 21422 3012
rect 21821 3009 21833 3012
rect 21867 3009 21879 3043
rect 21821 3003 21879 3009
rect 22088 3003 22100 3049
rect 22152 3040 22158 3052
rect 23937 3043 23995 3049
rect 22152 3012 22188 3040
rect 22094 3000 22100 3003
rect 22152 3000 22158 3012
rect 23937 3009 23949 3043
rect 23983 3040 23995 3043
rect 24136 3040 24164 3068
rect 24489 3043 24547 3049
rect 24489 3040 24501 3043
rect 23983 3012 24072 3040
rect 24136 3012 24501 3040
rect 23983 3009 23995 3012
rect 23937 3003 23995 3009
rect 23753 2907 23811 2913
rect 23753 2904 23765 2907
rect 15488 2876 20300 2904
rect 22756 2876 23765 2904
rect 16114 2836 16120 2848
rect 15212 2808 16120 2836
rect 16114 2796 16120 2808
rect 16172 2796 16178 2848
rect 18325 2839 18383 2845
rect 18325 2805 18337 2839
rect 18371 2836 18383 2839
rect 18598 2836 18604 2848
rect 18371 2808 18604 2836
rect 18371 2805 18383 2808
rect 18325 2799 18383 2805
rect 18598 2796 18604 2808
rect 18656 2836 18662 2848
rect 20162 2836 20168 2848
rect 18656 2808 20168 2836
rect 18656 2796 18662 2808
rect 20162 2796 20168 2808
rect 20220 2796 20226 2848
rect 20530 2796 20536 2848
rect 20588 2836 20594 2848
rect 20717 2839 20775 2845
rect 20717 2836 20729 2839
rect 20588 2808 20729 2836
rect 20588 2796 20594 2808
rect 20717 2805 20729 2808
rect 20763 2805 20775 2839
rect 20717 2799 20775 2805
rect 22186 2796 22192 2848
rect 22244 2836 22250 2848
rect 22756 2836 22784 2876
rect 23753 2873 23765 2876
rect 23799 2873 23811 2907
rect 23753 2867 23811 2873
rect 22244 2808 22784 2836
rect 24044 2836 24072 3012
rect 24489 3009 24501 3012
rect 24535 3009 24547 3043
rect 24489 3003 24547 3009
rect 24578 3000 24584 3052
rect 24636 3040 24642 3052
rect 24745 3043 24803 3049
rect 24745 3040 24757 3043
rect 24636 3012 24757 3040
rect 24636 3000 24642 3012
rect 24745 3009 24757 3012
rect 24791 3009 24803 3043
rect 24745 3003 24803 3009
rect 26436 2836 26464 3071
rect 27430 3068 27436 3080
rect 27488 3068 27494 3120
rect 28074 3068 28080 3120
rect 28132 3117 28138 3120
rect 28132 3108 28144 3117
rect 28132 3080 28177 3108
rect 28132 3071 28144 3080
rect 28132 3068 28138 3071
rect 29638 3068 29644 3120
rect 29696 3108 29702 3120
rect 29948 3111 30006 3117
rect 29948 3108 29960 3111
rect 29696 3080 29960 3108
rect 29696 3068 29702 3080
rect 29948 3077 29960 3080
rect 29994 3108 30006 3111
rect 30190 3108 30196 3120
rect 29994 3080 30196 3108
rect 29994 3077 30006 3080
rect 29948 3071 30006 3077
rect 30190 3068 30196 3080
rect 30248 3068 30254 3120
rect 32766 3108 32772 3120
rect 31404 3080 32772 3108
rect 28350 3040 28356 3052
rect 28311 3012 28356 3040
rect 28350 3000 28356 3012
rect 28408 3000 28414 3052
rect 30098 3000 30104 3052
rect 30156 3040 30162 3052
rect 30558 3040 30564 3052
rect 30156 3012 30564 3040
rect 30156 3000 30162 3012
rect 30558 3000 30564 3012
rect 30616 3040 30622 3052
rect 30653 3043 30711 3049
rect 30653 3040 30665 3043
rect 30616 3012 30665 3040
rect 30616 3000 30622 3012
rect 30653 3009 30665 3012
rect 30699 3009 30711 3043
rect 30653 3003 30711 3009
rect 31018 3000 31024 3052
rect 31076 3040 31082 3052
rect 31404 3049 31432 3080
rect 32766 3068 32772 3080
rect 32824 3068 32830 3120
rect 36204 3111 36262 3117
rect 36204 3077 36216 3111
rect 36250 3108 36262 3111
rect 37274 3108 37280 3120
rect 36250 3080 37280 3108
rect 36250 3077 36262 3080
rect 36204 3071 36262 3077
rect 37274 3068 37280 3080
rect 37332 3068 37338 3120
rect 37642 3068 37648 3120
rect 37700 3108 37706 3120
rect 38010 3108 38016 3120
rect 37700 3080 38016 3108
rect 37700 3068 37706 3080
rect 38010 3068 38016 3080
rect 38068 3068 38074 3120
rect 31389 3043 31447 3049
rect 31389 3040 31401 3043
rect 31076 3012 31401 3040
rect 31076 3000 31082 3012
rect 31389 3009 31401 3012
rect 31435 3009 31447 3043
rect 31389 3003 31447 3009
rect 31754 3000 31760 3052
rect 31812 3040 31818 3052
rect 32381 3043 32439 3049
rect 32381 3040 32393 3043
rect 31812 3012 32393 3040
rect 31812 3000 31818 3012
rect 32381 3009 32393 3012
rect 32427 3009 32439 3043
rect 34146 3040 34152 3052
rect 34107 3012 34152 3040
rect 32381 3003 32439 3009
rect 34146 3000 34152 3012
rect 34204 3000 34210 3052
rect 36354 3000 36360 3052
rect 36412 3040 36418 3052
rect 36449 3043 36507 3049
rect 36449 3040 36461 3043
rect 36412 3012 36461 3040
rect 36412 3000 36418 3012
rect 36449 3009 36461 3012
rect 36495 3009 36507 3043
rect 36449 3003 36507 3009
rect 30193 2975 30251 2981
rect 30193 2941 30205 2975
rect 30239 2972 30251 2975
rect 31478 2972 31484 2984
rect 30239 2944 31484 2972
rect 30239 2941 30251 2944
rect 30193 2935 30251 2941
rect 31478 2932 31484 2944
rect 31536 2972 31542 2984
rect 32122 2972 32128 2984
rect 31536 2944 32128 2972
rect 31536 2932 31542 2944
rect 32122 2932 32128 2944
rect 32180 2932 32186 2984
rect 26878 2864 26884 2916
rect 26936 2904 26942 2916
rect 26973 2907 27031 2913
rect 26973 2904 26985 2907
rect 26936 2876 26985 2904
rect 26936 2864 26942 2876
rect 26973 2873 26985 2876
rect 27019 2873 27031 2907
rect 31294 2904 31300 2916
rect 26973 2867 27031 2873
rect 30208 2876 31300 2904
rect 24044 2808 26464 2836
rect 22244 2796 22250 2808
rect 29454 2796 29460 2848
rect 29512 2836 29518 2848
rect 30208 2836 30236 2876
rect 31294 2864 31300 2876
rect 31352 2864 31358 2916
rect 34164 2904 34192 3000
rect 33060 2876 34192 2904
rect 29512 2808 30236 2836
rect 29512 2796 29518 2808
rect 30466 2796 30472 2848
rect 30524 2836 30530 2848
rect 33060 2836 33088 2876
rect 33502 2836 33508 2848
rect 30524 2808 33088 2836
rect 33463 2808 33508 2836
rect 30524 2796 30530 2808
rect 33502 2796 33508 2808
rect 33560 2796 33566 2848
rect 34330 2796 34336 2848
rect 34388 2836 34394 2848
rect 37550 2836 37556 2848
rect 34388 2808 37556 2836
rect 34388 2796 34394 2808
rect 37550 2796 37556 2808
rect 37608 2796 37614 2848
rect 37921 2839 37979 2845
rect 37921 2805 37933 2839
rect 37967 2836 37979 2839
rect 38286 2836 38292 2848
rect 37967 2808 38292 2836
rect 37967 2805 37979 2808
rect 37921 2799 37979 2805
rect 38286 2796 38292 2808
rect 38344 2796 38350 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 7745 2635 7803 2641
rect 7745 2601 7757 2635
rect 7791 2632 7803 2635
rect 8662 2632 8668 2644
rect 7791 2604 8668 2632
rect 7791 2601 7803 2604
rect 7745 2595 7803 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 9674 2632 9680 2644
rect 9048 2604 9680 2632
rect 7101 2567 7159 2573
rect 7101 2533 7113 2567
rect 7147 2564 7159 2567
rect 8389 2567 8447 2573
rect 7147 2536 8340 2564
rect 7147 2533 7159 2536
rect 7101 2527 7159 2533
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 7466 2496 7472 2508
rect 4111 2468 7472 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 7466 2456 7472 2468
rect 7524 2456 7530 2508
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 1762 2428 1768 2440
rect 1719 2400 1768 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 1762 2388 1768 2400
rect 1820 2388 1826 2440
rect 2314 2388 2320 2440
rect 2372 2428 2378 2440
rect 2409 2431 2467 2437
rect 2409 2428 2421 2431
rect 2372 2400 2421 2428
rect 2372 2388 2378 2400
rect 2409 2397 2421 2400
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 2700 2360 2728 2391
rect 2866 2388 2872 2440
rect 2924 2428 2930 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 2924 2400 3801 2428
rect 2924 2388 2930 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 5629 2431 5687 2437
rect 5629 2428 5641 2431
rect 5592 2400 5641 2428
rect 5592 2388 5598 2400
rect 5629 2397 5641 2400
rect 5675 2397 5687 2431
rect 5629 2391 5687 2397
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 7282 2428 7288 2440
rect 6963 2400 7288 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 8202 2428 8208 2440
rect 7607 2400 8064 2428
rect 8163 2400 8208 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 5718 2360 5724 2372
rect 2700 2332 5724 2360
rect 5718 2320 5724 2332
rect 5776 2320 5782 2372
rect 8036 2360 8064 2400
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 8312 2428 8340 2536
rect 8389 2533 8401 2567
rect 8435 2564 8447 2567
rect 9048 2564 9076 2604
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 9861 2635 9919 2641
rect 9861 2601 9873 2635
rect 9907 2632 9919 2635
rect 9950 2632 9956 2644
rect 9907 2604 9956 2632
rect 9907 2601 9919 2604
rect 9861 2595 9919 2601
rect 9950 2592 9956 2604
rect 10008 2592 10014 2644
rect 10689 2635 10747 2641
rect 10689 2601 10701 2635
rect 10735 2632 10747 2635
rect 11882 2632 11888 2644
rect 10735 2604 11888 2632
rect 10735 2601 10747 2604
rect 10689 2595 10747 2601
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12342 2592 12348 2644
rect 12400 2632 12406 2644
rect 14550 2632 14556 2644
rect 12400 2604 14556 2632
rect 12400 2592 12406 2604
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 14826 2632 14832 2644
rect 14787 2604 14832 2632
rect 14826 2592 14832 2604
rect 14884 2592 14890 2644
rect 16117 2635 16175 2641
rect 16117 2601 16129 2635
rect 16163 2632 16175 2635
rect 16850 2632 16856 2644
rect 16163 2604 16856 2632
rect 16163 2601 16175 2604
rect 16117 2595 16175 2601
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 17129 2635 17187 2641
rect 17129 2601 17141 2635
rect 17175 2632 17187 2635
rect 18322 2632 18328 2644
rect 17175 2604 18328 2632
rect 17175 2601 17187 2604
rect 17129 2595 17187 2601
rect 18322 2592 18328 2604
rect 18380 2592 18386 2644
rect 19426 2592 19432 2644
rect 19484 2632 19490 2644
rect 19981 2635 20039 2641
rect 19981 2632 19993 2635
rect 19484 2604 19993 2632
rect 19484 2592 19490 2604
rect 19981 2601 19993 2604
rect 20027 2601 20039 2635
rect 20438 2632 20444 2644
rect 20399 2604 20444 2632
rect 19981 2595 20039 2601
rect 20438 2592 20444 2604
rect 20496 2592 20502 2644
rect 26510 2632 26516 2644
rect 20548 2604 26516 2632
rect 8435 2536 9076 2564
rect 9217 2567 9275 2573
rect 8435 2533 8447 2536
rect 8389 2527 8447 2533
rect 9217 2533 9229 2567
rect 9263 2564 9275 2567
rect 11790 2564 11796 2576
rect 9263 2536 11796 2564
rect 9263 2533 9275 2536
rect 9217 2527 9275 2533
rect 11790 2524 11796 2536
rect 11848 2524 11854 2576
rect 12250 2524 12256 2576
rect 12308 2564 12314 2576
rect 20548 2564 20576 2604
rect 26510 2592 26516 2604
rect 26568 2592 26574 2644
rect 26602 2592 26608 2644
rect 26660 2632 26666 2644
rect 28537 2635 28595 2641
rect 28537 2632 28549 2635
rect 26660 2604 28549 2632
rect 26660 2592 26666 2604
rect 28537 2601 28549 2604
rect 28583 2601 28595 2635
rect 28537 2595 28595 2601
rect 30650 2592 30656 2644
rect 30708 2632 30714 2644
rect 30837 2635 30895 2641
rect 30837 2632 30849 2635
rect 30708 2604 30849 2632
rect 30708 2592 30714 2604
rect 30837 2601 30849 2604
rect 30883 2601 30895 2635
rect 30837 2595 30895 2601
rect 31662 2592 31668 2644
rect 31720 2632 31726 2644
rect 31720 2604 33548 2632
rect 31720 2592 31726 2604
rect 22281 2567 22339 2573
rect 22281 2564 22293 2567
rect 12308 2536 20576 2564
rect 22066 2536 22293 2564
rect 12308 2524 12314 2536
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2496 10379 2499
rect 11054 2496 11060 2508
rect 10367 2468 11060 2496
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 11256 2468 13400 2496
rect 8478 2428 8484 2440
rect 8312 2400 8484 2428
rect 8478 2388 8484 2400
rect 8536 2388 8542 2440
rect 9030 2428 9036 2440
rect 8991 2400 9036 2428
rect 9030 2388 9036 2400
rect 9088 2388 9094 2440
rect 9490 2388 9496 2440
rect 9548 2428 9554 2440
rect 9677 2431 9735 2437
rect 9677 2428 9689 2431
rect 9548 2400 9689 2428
rect 9548 2388 9554 2400
rect 9677 2397 9689 2400
rect 9723 2397 9735 2431
rect 10502 2428 10508 2440
rect 10463 2400 10508 2428
rect 9677 2391 9735 2397
rect 8294 2360 8300 2372
rect 8036 2332 8300 2360
rect 8294 2320 8300 2332
rect 8352 2320 8358 2372
rect 9692 2360 9720 2391
rect 10502 2388 10508 2400
rect 10560 2388 10566 2440
rect 11146 2360 11152 2372
rect 9692 2332 11152 2360
rect 11146 2320 11152 2332
rect 11204 2320 11210 2372
rect 1854 2292 1860 2304
rect 1815 2264 1860 2292
rect 1854 2252 1860 2264
rect 1912 2252 1918 2304
rect 5166 2292 5172 2304
rect 5127 2264 5172 2292
rect 5166 2252 5172 2264
rect 5224 2252 5230 2304
rect 5810 2292 5816 2304
rect 5771 2264 5816 2292
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 6457 2295 6515 2301
rect 6457 2261 6469 2295
rect 6503 2292 6515 2295
rect 11256 2292 11284 2468
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12434 2428 12440 2440
rect 12115 2400 12440 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 12618 2388 12624 2440
rect 12676 2428 12682 2440
rect 13372 2437 13400 2468
rect 13446 2456 13452 2508
rect 13504 2496 13510 2508
rect 13504 2468 14688 2496
rect 13504 2456 13510 2468
rect 14660 2437 14688 2468
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 17218 2496 17224 2508
rect 15252 2468 17224 2496
rect 15252 2456 15258 2468
rect 15304 2437 15332 2468
rect 17218 2456 17224 2468
rect 17276 2456 17282 2508
rect 19150 2496 19156 2508
rect 17696 2468 19156 2496
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 12676 2400 12725 2428
rect 12676 2388 12682 2400
rect 12713 2397 12725 2400
rect 12759 2397 12771 2431
rect 12713 2391 12771 2397
rect 13357 2431 13415 2437
rect 13357 2397 13369 2431
rect 13403 2428 13415 2431
rect 14645 2431 14703 2437
rect 13403 2400 14596 2428
rect 13403 2397 13415 2400
rect 13357 2391 13415 2397
rect 14458 2360 14464 2372
rect 12912 2332 14464 2360
rect 11606 2292 11612 2304
rect 6503 2264 11284 2292
rect 11567 2264 11612 2292
rect 6503 2261 6515 2264
rect 6457 2255 6515 2261
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 12253 2295 12311 2301
rect 12253 2261 12265 2295
rect 12299 2292 12311 2295
rect 12342 2292 12348 2304
rect 12299 2264 12348 2292
rect 12299 2261 12311 2264
rect 12253 2255 12311 2261
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 12912 2301 12940 2332
rect 14458 2320 14464 2332
rect 14516 2320 14522 2372
rect 14568 2360 14596 2400
rect 14645 2397 14657 2431
rect 14691 2428 14703 2431
rect 15289 2431 15347 2437
rect 14691 2400 15148 2428
rect 14691 2397 14703 2400
rect 14645 2391 14703 2397
rect 15010 2360 15016 2372
rect 14568 2332 15016 2360
rect 15010 2320 15016 2332
rect 15068 2320 15074 2372
rect 15120 2360 15148 2400
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 16666 2428 16672 2440
rect 15335 2400 15369 2428
rect 15488 2400 16672 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15488 2360 15516 2400
rect 16666 2388 16672 2400
rect 16724 2388 16730 2440
rect 16942 2428 16948 2440
rect 16903 2400 16948 2428
rect 16942 2388 16948 2400
rect 17000 2388 17006 2440
rect 17696 2437 17724 2468
rect 19150 2456 19156 2468
rect 19208 2456 19214 2508
rect 19334 2496 19340 2508
rect 19295 2468 19340 2496
rect 19334 2456 19340 2468
rect 19392 2456 19398 2508
rect 20162 2456 20168 2508
rect 20220 2496 20226 2508
rect 22066 2496 22094 2536
rect 22281 2533 22293 2536
rect 22327 2533 22339 2567
rect 22281 2527 22339 2533
rect 24394 2524 24400 2576
rect 24452 2564 24458 2576
rect 25961 2567 26019 2573
rect 25961 2564 25973 2567
rect 24452 2536 25973 2564
rect 24452 2524 24458 2536
rect 25961 2533 25973 2536
rect 26007 2533 26019 2567
rect 27065 2567 27123 2573
rect 27065 2564 27077 2567
rect 25961 2527 26019 2533
rect 26068 2536 27077 2564
rect 20220 2468 22094 2496
rect 23661 2499 23719 2505
rect 20220 2456 20226 2468
rect 23661 2465 23673 2499
rect 23707 2496 23719 2499
rect 24118 2496 24124 2508
rect 23707 2468 24124 2496
rect 23707 2465 23719 2468
rect 23661 2459 23719 2465
rect 24118 2456 24124 2468
rect 24176 2456 24182 2508
rect 25498 2456 25504 2508
rect 25556 2496 25562 2508
rect 26068 2496 26096 2536
rect 27065 2533 27077 2536
rect 27111 2533 27123 2567
rect 28994 2564 29000 2576
rect 27065 2527 27123 2533
rect 27172 2536 29000 2564
rect 27172 2496 27200 2536
rect 28994 2524 29000 2536
rect 29052 2524 29058 2576
rect 30377 2567 30435 2573
rect 30377 2533 30389 2567
rect 30423 2564 30435 2567
rect 32490 2564 32496 2576
rect 30423 2536 32496 2564
rect 30423 2533 30435 2536
rect 30377 2527 30435 2533
rect 32490 2524 32496 2536
rect 32548 2524 32554 2576
rect 33520 2564 33548 2604
rect 33594 2592 33600 2644
rect 33652 2632 33658 2644
rect 33965 2635 34023 2641
rect 33965 2632 33977 2635
rect 33652 2604 33977 2632
rect 33652 2592 33658 2604
rect 33965 2601 33977 2604
rect 34011 2601 34023 2635
rect 33965 2595 34023 2601
rect 36446 2592 36452 2644
rect 36504 2632 36510 2644
rect 36504 2604 36768 2632
rect 36504 2592 36510 2604
rect 35345 2567 35403 2573
rect 35345 2564 35357 2567
rect 33520 2536 35357 2564
rect 35345 2533 35357 2536
rect 35391 2533 35403 2567
rect 35345 2527 35403 2533
rect 25556 2468 26096 2496
rect 26160 2468 27200 2496
rect 27908 2468 31616 2496
rect 25556 2456 25562 2468
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2397 17739 2431
rect 17954 2428 17960 2440
rect 17681 2391 17739 2397
rect 17788 2400 17960 2428
rect 15120 2332 15516 2360
rect 12897 2295 12955 2301
rect 12897 2261 12909 2295
rect 12943 2261 12955 2295
rect 13538 2292 13544 2304
rect 13499 2264 13544 2292
rect 12897 2255 12955 2261
rect 13538 2252 13544 2264
rect 13596 2252 13602 2304
rect 14182 2292 14188 2304
rect 14143 2264 14188 2292
rect 14182 2252 14188 2264
rect 14240 2252 14246 2304
rect 15473 2295 15531 2301
rect 15473 2261 15485 2295
rect 15519 2292 15531 2295
rect 17788 2292 17816 2400
rect 17954 2388 17960 2400
rect 18012 2388 18018 2440
rect 18414 2428 18420 2440
rect 18375 2400 18420 2428
rect 18414 2388 18420 2400
rect 18472 2428 18478 2440
rect 18690 2428 18696 2440
rect 18472 2400 18696 2428
rect 18472 2388 18478 2400
rect 18690 2388 18696 2400
rect 18748 2388 18754 2440
rect 19521 2431 19579 2437
rect 19521 2397 19533 2431
rect 19567 2428 19579 2431
rect 20714 2428 20720 2440
rect 19567 2400 20720 2428
rect 19567 2397 19579 2400
rect 19521 2391 19579 2397
rect 20714 2388 20720 2400
rect 20772 2388 20778 2440
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 22462 2428 22468 2440
rect 21315 2400 22468 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 22462 2388 22468 2400
rect 22520 2388 22526 2440
rect 24673 2431 24731 2437
rect 24673 2397 24685 2431
rect 24719 2428 24731 2431
rect 25038 2428 25044 2440
rect 24719 2400 25044 2428
rect 24719 2397 24731 2400
rect 24673 2391 24731 2397
rect 25038 2388 25044 2400
rect 25096 2388 25102 2440
rect 26160 2437 26188 2468
rect 25409 2431 25467 2437
rect 25409 2397 25421 2431
rect 25455 2397 25467 2431
rect 25409 2391 25467 2397
rect 26145 2431 26203 2437
rect 26145 2397 26157 2431
rect 26191 2397 26203 2431
rect 26326 2428 26332 2440
rect 26145 2391 26203 2397
rect 26252 2400 26332 2428
rect 18874 2360 18880 2372
rect 17880 2332 18880 2360
rect 17880 2301 17908 2332
rect 18874 2320 18880 2332
rect 18932 2320 18938 2372
rect 19610 2360 19616 2372
rect 19571 2332 19616 2360
rect 19610 2320 19616 2332
rect 19668 2320 19674 2372
rect 20070 2320 20076 2372
rect 20128 2360 20134 2372
rect 23394 2363 23452 2369
rect 23394 2360 23406 2363
rect 20128 2332 23406 2360
rect 20128 2320 20134 2332
rect 23394 2329 23406 2332
rect 23440 2329 23452 2363
rect 25424 2360 25452 2391
rect 26252 2360 26280 2400
rect 26326 2388 26332 2400
rect 26384 2388 26390 2440
rect 27249 2431 27307 2437
rect 27249 2397 27261 2431
rect 27295 2424 27307 2431
rect 27908 2428 27936 2468
rect 27356 2424 27936 2428
rect 27295 2400 27936 2424
rect 27985 2431 28043 2437
rect 27295 2397 27384 2400
rect 27249 2396 27384 2397
rect 27985 2397 27997 2431
rect 28031 2397 28043 2431
rect 28718 2428 28724 2440
rect 28679 2400 28724 2428
rect 27249 2391 27307 2396
rect 27985 2391 28043 2397
rect 23394 2323 23452 2329
rect 23492 2332 25268 2360
rect 25424 2332 26280 2360
rect 26344 2332 27844 2360
rect 15519 2264 17816 2292
rect 17865 2295 17923 2301
rect 15519 2261 15531 2264
rect 15473 2255 15531 2261
rect 17865 2261 17877 2295
rect 17911 2261 17923 2295
rect 17865 2255 17923 2261
rect 17954 2252 17960 2304
rect 18012 2292 18018 2304
rect 18506 2292 18512 2304
rect 18012 2264 18512 2292
rect 18012 2252 18018 2264
rect 18506 2252 18512 2264
rect 18564 2252 18570 2304
rect 18601 2295 18659 2301
rect 18601 2261 18613 2295
rect 18647 2292 18659 2295
rect 19426 2292 19432 2304
rect 18647 2264 19432 2292
rect 18647 2261 18659 2264
rect 18601 2255 18659 2261
rect 19426 2252 19432 2264
rect 19484 2252 19490 2304
rect 21082 2292 21088 2304
rect 21043 2264 21088 2292
rect 21082 2252 21088 2264
rect 21140 2252 21146 2304
rect 23290 2252 23296 2304
rect 23348 2292 23354 2304
rect 23492 2292 23520 2332
rect 24486 2292 24492 2304
rect 23348 2264 23520 2292
rect 24447 2264 24492 2292
rect 23348 2252 23354 2264
rect 24486 2252 24492 2264
rect 24544 2252 24550 2304
rect 25240 2301 25268 2332
rect 25225 2295 25283 2301
rect 25225 2261 25237 2295
rect 25271 2261 25283 2295
rect 25225 2255 25283 2261
rect 26050 2252 26056 2304
rect 26108 2292 26114 2304
rect 26344 2292 26372 2332
rect 27816 2301 27844 2332
rect 26108 2264 26372 2292
rect 27801 2295 27859 2301
rect 26108 2252 26114 2264
rect 27801 2261 27813 2295
rect 27847 2261 27859 2295
rect 28000 2292 28028 2391
rect 28718 2388 28724 2400
rect 28776 2388 28782 2440
rect 29362 2428 29368 2440
rect 28828 2400 29368 2428
rect 28074 2320 28080 2372
rect 28132 2360 28138 2372
rect 28828 2360 28856 2400
rect 29362 2388 29368 2400
rect 29420 2428 29426 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29420 2400 29745 2428
rect 29420 2388 29426 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30193 2431 30251 2437
rect 30193 2397 30205 2431
rect 30239 2397 30251 2431
rect 30193 2391 30251 2397
rect 31021 2431 31079 2437
rect 31021 2397 31033 2431
rect 31067 2428 31079 2431
rect 31294 2428 31300 2440
rect 31067 2400 31300 2428
rect 31067 2397 31079 2400
rect 31021 2391 31079 2397
rect 28132 2332 28856 2360
rect 28132 2320 28138 2332
rect 28994 2320 29000 2372
rect 29052 2360 29058 2372
rect 29822 2360 29828 2372
rect 29052 2332 29828 2360
rect 29052 2320 29058 2332
rect 29822 2320 29828 2332
rect 29880 2360 29886 2372
rect 30208 2360 30236 2391
rect 31294 2388 31300 2400
rect 31352 2388 31358 2440
rect 31588 2437 31616 2468
rect 32122 2456 32128 2508
rect 32180 2496 32186 2508
rect 36740 2505 36768 2604
rect 32585 2499 32643 2505
rect 32585 2496 32597 2499
rect 32180 2468 32597 2496
rect 32180 2456 32186 2468
rect 32585 2465 32597 2468
rect 32631 2465 32643 2499
rect 32585 2459 32643 2465
rect 36725 2499 36783 2505
rect 36725 2465 36737 2499
rect 36771 2465 36783 2499
rect 37550 2496 37556 2508
rect 37511 2468 37556 2496
rect 36725 2459 36783 2465
rect 37550 2456 37556 2468
rect 37608 2456 37614 2508
rect 31573 2431 31631 2437
rect 31573 2397 31585 2431
rect 31619 2428 31631 2431
rect 34238 2428 34244 2440
rect 31619 2400 34244 2428
rect 31619 2397 31631 2400
rect 31573 2391 31631 2397
rect 34238 2388 34244 2400
rect 34296 2388 34302 2440
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34848 2400 34897 2428
rect 34848 2388 34854 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 36469 2431 36527 2437
rect 36469 2397 36481 2431
rect 36515 2428 36527 2431
rect 36630 2428 36636 2440
rect 36515 2400 36636 2428
rect 36515 2397 36527 2400
rect 36469 2391 36527 2397
rect 36630 2388 36636 2400
rect 36688 2388 36694 2440
rect 37090 2388 37096 2440
rect 37148 2428 37154 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 37148 2400 37289 2428
rect 37148 2388 37154 2400
rect 37277 2397 37289 2400
rect 37323 2428 37335 2431
rect 37826 2428 37832 2440
rect 37323 2400 37832 2428
rect 37323 2397 37335 2400
rect 37277 2391 37335 2397
rect 37826 2388 37832 2400
rect 37884 2388 37890 2440
rect 29880 2332 30236 2360
rect 32852 2363 32910 2369
rect 29880 2320 29886 2332
rect 32852 2329 32864 2363
rect 32898 2360 32910 2363
rect 32898 2332 34744 2360
rect 32898 2329 32910 2332
rect 32852 2323 32910 2329
rect 29086 2292 29092 2304
rect 28000 2264 29092 2292
rect 27801 2255 27859 2261
rect 29086 2252 29092 2264
rect 29144 2252 29150 2304
rect 29546 2292 29552 2304
rect 29507 2264 29552 2292
rect 29546 2252 29552 2264
rect 29604 2252 29610 2304
rect 34716 2301 34744 2332
rect 34701 2295 34759 2301
rect 34701 2261 34713 2295
rect 34747 2261 34759 2295
rect 34701 2255 34759 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 1854 2048 1860 2100
rect 1912 2088 1918 2100
rect 1912 2060 2774 2088
rect 1912 2048 1918 2060
rect 2746 2020 2774 2060
rect 5810 2048 5816 2100
rect 5868 2088 5874 2100
rect 9858 2088 9864 2100
rect 5868 2060 9864 2088
rect 5868 2048 5874 2060
rect 9858 2048 9864 2060
rect 9916 2048 9922 2100
rect 10962 2048 10968 2100
rect 11020 2088 11026 2100
rect 13446 2088 13452 2100
rect 11020 2060 13452 2088
rect 11020 2048 11026 2060
rect 13446 2048 13452 2060
rect 13504 2048 13510 2100
rect 13538 2048 13544 2100
rect 13596 2088 13602 2100
rect 16574 2088 16580 2100
rect 13596 2060 16580 2088
rect 13596 2048 13602 2060
rect 16574 2048 16580 2060
rect 16632 2048 16638 2100
rect 21634 2048 21640 2100
rect 21692 2088 21698 2100
rect 24486 2088 24492 2100
rect 21692 2060 24492 2088
rect 21692 2048 21698 2060
rect 24486 2048 24492 2060
rect 24544 2048 24550 2100
rect 26510 2048 26516 2100
rect 26568 2088 26574 2100
rect 29638 2088 29644 2100
rect 26568 2060 29644 2088
rect 26568 2048 26574 2060
rect 29638 2048 29644 2060
rect 29696 2048 29702 2100
rect 8754 2020 8760 2032
rect 2746 1992 8760 2020
rect 8754 1980 8760 1992
rect 8812 1980 8818 2032
rect 14182 1980 14188 2032
rect 14240 2020 14246 2032
rect 18414 2020 18420 2032
rect 14240 1992 18420 2020
rect 14240 1980 14246 1992
rect 18414 1980 18420 1992
rect 18472 1980 18478 2032
rect 5718 1912 5724 1964
rect 5776 1952 5782 1964
rect 8570 1952 8576 1964
rect 5776 1924 8576 1952
rect 5776 1912 5782 1924
rect 8570 1912 8576 1924
rect 8628 1912 8634 1964
rect 17862 1912 17868 1964
rect 17920 1952 17926 1964
rect 29546 1952 29552 1964
rect 17920 1924 29552 1952
rect 17920 1912 17926 1924
rect 29546 1912 29552 1924
rect 29604 1912 29610 1964
rect 5166 1844 5172 1896
rect 5224 1884 5230 1896
rect 12434 1884 12440 1896
rect 5224 1856 12440 1884
rect 5224 1844 5230 1856
rect 12434 1844 12440 1856
rect 12492 1884 12498 1896
rect 13354 1884 13360 1896
rect 12492 1856 13360 1884
rect 12492 1844 12498 1856
rect 13354 1844 13360 1856
rect 13412 1844 13418 1896
rect 13722 1844 13728 1896
rect 13780 1884 13786 1896
rect 20070 1884 20076 1896
rect 13780 1856 20076 1884
rect 13780 1844 13786 1856
rect 20070 1844 20076 1856
rect 20128 1844 20134 1896
rect 11606 1776 11612 1828
rect 11664 1816 11670 1828
rect 16942 1816 16948 1828
rect 11664 1788 16948 1816
rect 11664 1776 11670 1788
rect 16942 1776 16948 1788
rect 17000 1776 17006 1828
rect 5534 1708 5540 1760
rect 5592 1748 5598 1760
rect 6178 1748 6184 1760
rect 5592 1720 6184 1748
rect 5592 1708 5598 1720
rect 6178 1708 6184 1720
rect 6236 1708 6242 1760
rect 8202 1708 8208 1760
rect 8260 1748 8266 1760
rect 9490 1748 9496 1760
rect 8260 1720 9496 1748
rect 8260 1708 8266 1720
rect 9490 1708 9496 1720
rect 9548 1708 9554 1760
rect 12618 1708 12624 1760
rect 12676 1748 12682 1760
rect 14458 1748 14464 1760
rect 12676 1720 14464 1748
rect 12676 1708 12682 1720
rect 14458 1708 14464 1720
rect 14516 1708 14522 1760
rect 16850 1368 16856 1420
rect 16908 1408 16914 1420
rect 17770 1408 17776 1420
rect 16908 1380 17776 1408
rect 16908 1368 16914 1380
rect 17770 1368 17776 1380
rect 17828 1368 17834 1420
<< via1 >>
rect 21272 37680 21324 37732
rect 23848 37680 23900 37732
rect 13452 37612 13504 37664
rect 26240 37612 26292 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 23848 37451 23900 37460
rect 9956 37340 10008 37392
rect 23848 37417 23857 37451
rect 23857 37417 23891 37451
rect 23891 37417 23900 37451
rect 23848 37408 23900 37417
rect 28448 37408 28500 37460
rect 29368 37408 29420 37460
rect 35072 37340 35124 37392
rect 17776 37272 17828 37324
rect 1768 37204 1820 37256
rect 2504 37247 2556 37256
rect 2504 37213 2513 37247
rect 2513 37213 2547 37247
rect 2547 37213 2556 37247
rect 2504 37204 2556 37213
rect 3240 37247 3292 37256
rect 3240 37213 3249 37247
rect 3249 37213 3283 37247
rect 3283 37213 3292 37247
rect 3240 37204 3292 37213
rect 4712 37204 4764 37256
rect 5816 37247 5868 37256
rect 5816 37213 5825 37247
rect 5825 37213 5859 37247
rect 5859 37213 5868 37247
rect 5816 37204 5868 37213
rect 7012 37136 7064 37188
rect 7380 37204 7432 37256
rect 8576 37204 8628 37256
rect 8300 37136 8352 37188
rect 2320 37111 2372 37120
rect 2320 37077 2329 37111
rect 2329 37077 2363 37111
rect 2363 37077 2372 37111
rect 2320 37068 2372 37077
rect 2872 37068 2924 37120
rect 4160 37111 4212 37120
rect 4160 37077 4169 37111
rect 4169 37077 4203 37111
rect 4203 37077 4212 37111
rect 4160 37068 4212 37077
rect 5080 37068 5132 37120
rect 5632 37111 5684 37120
rect 5632 37077 5641 37111
rect 5641 37077 5675 37111
rect 5675 37077 5684 37111
rect 5632 37068 5684 37077
rect 6736 37111 6788 37120
rect 6736 37077 6745 37111
rect 6745 37077 6779 37111
rect 6779 37077 6788 37111
rect 6736 37068 6788 37077
rect 7288 37068 7340 37120
rect 8392 37068 8444 37120
rect 9496 37068 9548 37120
rect 10048 37111 10100 37120
rect 10048 37077 10057 37111
rect 10057 37077 10091 37111
rect 10091 37077 10100 37111
rect 10048 37068 10100 37077
rect 10324 37204 10376 37256
rect 12072 37247 12124 37256
rect 12072 37213 12081 37247
rect 12081 37213 12115 37247
rect 12115 37213 12124 37247
rect 12072 37204 12124 37213
rect 12532 37247 12584 37256
rect 12532 37213 12541 37247
rect 12541 37213 12575 37247
rect 12575 37213 12584 37247
rect 12532 37204 12584 37213
rect 13544 37247 13596 37256
rect 13544 37213 13553 37247
rect 13553 37213 13587 37247
rect 13587 37213 13596 37247
rect 13544 37204 13596 37213
rect 14648 37247 14700 37256
rect 14648 37213 14657 37247
rect 14657 37213 14691 37247
rect 14691 37213 14700 37247
rect 14648 37204 14700 37213
rect 15384 37247 15436 37256
rect 15384 37213 15393 37247
rect 15393 37213 15427 37247
rect 15427 37213 15436 37247
rect 15384 37204 15436 37213
rect 15844 37247 15896 37256
rect 15844 37213 15853 37247
rect 15853 37213 15887 37247
rect 15887 37213 15896 37247
rect 15844 37204 15896 37213
rect 17684 37204 17736 37256
rect 10416 37136 10468 37188
rect 11060 37136 11112 37188
rect 16856 37136 16908 37188
rect 19340 37204 19392 37256
rect 19984 37204 20036 37256
rect 20168 37204 20220 37256
rect 20444 37204 20496 37256
rect 21180 37204 21232 37256
rect 34244 37272 34296 37324
rect 22100 37204 22152 37256
rect 23296 37247 23348 37256
rect 20812 37136 20864 37188
rect 11152 37068 11204 37120
rect 11704 37068 11756 37120
rect 12808 37068 12860 37120
rect 13360 37111 13412 37120
rect 13360 37077 13369 37111
rect 13369 37077 13403 37111
rect 13403 37077 13412 37111
rect 13360 37068 13412 37077
rect 14464 37111 14516 37120
rect 14464 37077 14473 37111
rect 14473 37077 14507 37111
rect 14507 37077 14516 37111
rect 14464 37068 14516 37077
rect 15200 37111 15252 37120
rect 15200 37077 15209 37111
rect 15209 37077 15243 37111
rect 15243 37077 15252 37111
rect 15200 37068 15252 37077
rect 16120 37068 16172 37120
rect 17224 37111 17276 37120
rect 17224 37077 17233 37111
rect 17233 37077 17267 37111
rect 17267 37077 17276 37111
rect 17224 37068 17276 37077
rect 20352 37068 20404 37120
rect 20904 37111 20956 37120
rect 20904 37077 20913 37111
rect 20913 37077 20947 37111
rect 20947 37077 20956 37111
rect 20904 37068 20956 37077
rect 20996 37068 21048 37120
rect 22192 37136 22244 37188
rect 23296 37213 23305 37247
rect 23305 37213 23339 37247
rect 23339 37213 23348 37247
rect 23296 37204 23348 37213
rect 23664 37204 23716 37256
rect 23388 37136 23440 37188
rect 25136 37204 25188 37256
rect 23112 37111 23164 37120
rect 23112 37077 23121 37111
rect 23121 37077 23155 37111
rect 23155 37077 23164 37111
rect 23112 37068 23164 37077
rect 24676 37068 24728 37120
rect 25044 37111 25096 37120
rect 25044 37077 25053 37111
rect 25053 37077 25087 37111
rect 25087 37077 25096 37111
rect 25044 37068 25096 37077
rect 25136 37068 25188 37120
rect 25320 37204 25372 37256
rect 27436 37204 27488 37256
rect 28080 37204 28132 37256
rect 29276 37204 29328 37256
rect 30380 37204 30432 37256
rect 31116 37204 31168 37256
rect 32220 37204 32272 37256
rect 32404 37247 32456 37256
rect 32404 37213 32413 37247
rect 32413 37213 32447 37247
rect 32447 37213 32456 37247
rect 32404 37204 32456 37213
rect 32496 37204 32548 37256
rect 30104 37136 30156 37188
rect 31576 37136 31628 37188
rect 34980 37204 35032 37256
rect 36084 37204 36136 37256
rect 25320 37068 25372 37120
rect 27160 37068 27212 37120
rect 27712 37068 27764 37120
rect 28264 37068 28316 37120
rect 29000 37068 29052 37120
rect 29920 37068 29972 37120
rect 31392 37068 31444 37120
rect 34796 37136 34848 37188
rect 35624 37179 35676 37188
rect 35624 37145 35658 37179
rect 35658 37145 35676 37179
rect 35624 37136 35676 37145
rect 35348 37068 35400 37120
rect 36728 37111 36780 37120
rect 36728 37077 36737 37111
rect 36737 37077 36771 37111
rect 36771 37077 36780 37111
rect 36728 37068 36780 37077
rect 38292 37068 38344 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 1768 36864 1820 36916
rect 3240 36864 3292 36916
rect 3424 36796 3476 36848
rect 4620 36864 4672 36916
rect 6184 36864 6236 36916
rect 7840 36864 7892 36916
rect 8944 36864 8996 36916
rect 10600 36864 10652 36916
rect 12440 36907 12492 36916
rect 12440 36873 12449 36907
rect 12449 36873 12483 36907
rect 12483 36873 12492 36907
rect 12440 36864 12492 36873
rect 13912 36864 13964 36916
rect 15568 36864 15620 36916
rect 16672 36864 16724 36916
rect 19432 36864 19484 36916
rect 19984 36907 20036 36916
rect 19984 36873 19993 36907
rect 19993 36873 20027 36907
rect 20027 36873 20036 36907
rect 19984 36864 20036 36873
rect 20812 36907 20864 36916
rect 20812 36873 20821 36907
rect 20821 36873 20855 36907
rect 20855 36873 20864 36907
rect 20812 36864 20864 36873
rect 21180 36864 21232 36916
rect 23664 36907 23716 36916
rect 9680 36796 9732 36848
rect 14648 36796 14700 36848
rect 18604 36796 18656 36848
rect 20996 36796 21048 36848
rect 5080 36728 5132 36780
rect 6644 36771 6696 36780
rect 6644 36737 6653 36771
rect 6653 36737 6687 36771
rect 6687 36737 6696 36771
rect 6644 36728 6696 36737
rect 8208 36771 8260 36780
rect 8208 36737 8217 36771
rect 8217 36737 8251 36771
rect 8251 36737 8260 36771
rect 8208 36728 8260 36737
rect 9312 36771 9364 36780
rect 9312 36737 9321 36771
rect 9321 36737 9355 36771
rect 9355 36737 9364 36771
rect 9312 36728 9364 36737
rect 10968 36771 11020 36780
rect 10968 36737 10977 36771
rect 10977 36737 11011 36771
rect 11011 36737 11020 36771
rect 10968 36728 11020 36737
rect 12624 36771 12676 36780
rect 12624 36737 12633 36771
rect 12633 36737 12667 36771
rect 12667 36737 12676 36771
rect 12624 36728 12676 36737
rect 14280 36771 14332 36780
rect 14280 36737 14289 36771
rect 14289 36737 14323 36771
rect 14323 36737 14332 36771
rect 14280 36728 14332 36737
rect 16028 36728 16080 36780
rect 17040 36771 17092 36780
rect 17040 36737 17049 36771
rect 17049 36737 17083 36771
rect 17083 36737 17092 36771
rect 17040 36728 17092 36737
rect 17868 36728 17920 36780
rect 6828 36592 6880 36644
rect 23664 36873 23673 36907
rect 23673 36873 23707 36907
rect 23707 36873 23716 36907
rect 23664 36864 23716 36873
rect 25412 36864 25464 36916
rect 24216 36796 24268 36848
rect 24768 36796 24820 36848
rect 28172 36864 28224 36916
rect 19432 36703 19484 36712
rect 19432 36669 19441 36703
rect 19441 36669 19475 36703
rect 19475 36669 19484 36703
rect 19432 36660 19484 36669
rect 21548 36660 21600 36712
rect 20260 36592 20312 36644
rect 23388 36728 23440 36780
rect 23020 36703 23072 36712
rect 23020 36669 23029 36703
rect 23029 36669 23063 36703
rect 23063 36669 23072 36703
rect 23020 36660 23072 36669
rect 23480 36660 23532 36712
rect 23388 36592 23440 36644
rect 5816 36567 5868 36576
rect 5816 36533 5825 36567
rect 5825 36533 5859 36567
rect 5859 36533 5868 36567
rect 5816 36524 5868 36533
rect 7380 36567 7432 36576
rect 7380 36533 7389 36567
rect 7389 36533 7423 36567
rect 7423 36533 7432 36567
rect 7380 36524 7432 36533
rect 10232 36567 10284 36576
rect 10232 36533 10241 36567
rect 10241 36533 10275 36567
rect 10275 36533 10284 36567
rect 10232 36524 10284 36533
rect 12532 36524 12584 36576
rect 17868 36524 17920 36576
rect 30472 36864 30524 36916
rect 34520 36864 34572 36916
rect 35072 36839 35124 36848
rect 35072 36805 35090 36839
rect 35090 36805 35124 36839
rect 35072 36796 35124 36805
rect 25504 36703 25556 36712
rect 25504 36669 25513 36703
rect 25513 36669 25547 36703
rect 25547 36669 25556 36703
rect 25504 36660 25556 36669
rect 29000 36660 29052 36712
rect 23756 36524 23808 36576
rect 26332 36592 26384 36644
rect 25964 36567 26016 36576
rect 25964 36533 25973 36567
rect 25973 36533 26007 36567
rect 26007 36533 26016 36567
rect 25964 36524 26016 36533
rect 26976 36567 27028 36576
rect 26976 36533 26985 36567
rect 26985 36533 27019 36567
rect 27019 36533 27028 36567
rect 26976 36524 27028 36533
rect 28448 36592 28500 36644
rect 30196 36703 30248 36712
rect 30196 36669 30205 36703
rect 30205 36669 30239 36703
rect 30239 36669 30248 36703
rect 30196 36660 30248 36669
rect 31300 36728 31352 36780
rect 35900 36728 35952 36780
rect 36452 36728 36504 36780
rect 38108 36728 38160 36780
rect 33784 36660 33836 36712
rect 35440 36592 35492 36644
rect 35900 36592 35952 36644
rect 36084 36592 36136 36644
rect 29276 36524 29328 36576
rect 33968 36567 34020 36576
rect 33968 36533 33977 36567
rect 33977 36533 34011 36567
rect 34011 36533 34020 36567
rect 33968 36524 34020 36533
rect 34980 36524 35032 36576
rect 37924 36524 37976 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 14280 36320 14332 36372
rect 16580 36320 16632 36372
rect 17776 36320 17828 36372
rect 19432 36363 19484 36372
rect 19432 36329 19441 36363
rect 19441 36329 19475 36363
rect 19475 36329 19484 36363
rect 19432 36320 19484 36329
rect 20168 36363 20220 36372
rect 20168 36329 20177 36363
rect 20177 36329 20211 36363
rect 20211 36329 20220 36363
rect 20168 36320 20220 36329
rect 6644 36252 6696 36304
rect 10048 36252 10100 36304
rect 17684 36252 17736 36304
rect 20076 36252 20128 36304
rect 2504 36184 2556 36236
rect 8760 36184 8812 36236
rect 9312 36184 9364 36236
rect 12716 36184 12768 36236
rect 15384 36184 15436 36236
rect 18420 36184 18472 36236
rect 8300 36116 8352 36168
rect 8944 36116 8996 36168
rect 10416 36159 10468 36168
rect 10416 36125 10425 36159
rect 10425 36125 10459 36159
rect 10459 36125 10468 36159
rect 10416 36116 10468 36125
rect 13176 36116 13228 36168
rect 13544 36159 13596 36168
rect 13544 36125 13553 36159
rect 13553 36125 13587 36159
rect 13587 36125 13596 36159
rect 13544 36116 13596 36125
rect 15752 36116 15804 36168
rect 18880 36116 18932 36168
rect 20628 36184 20680 36236
rect 21548 36227 21600 36236
rect 21548 36193 21557 36227
rect 21557 36193 21591 36227
rect 21591 36193 21600 36227
rect 21548 36184 21600 36193
rect 23112 36184 23164 36236
rect 7012 36048 7064 36100
rect 7564 36048 7616 36100
rect 10968 36048 11020 36100
rect 13636 36048 13688 36100
rect 20444 36048 20496 36100
rect 22376 36116 22428 36168
rect 22560 36159 22612 36168
rect 22560 36125 22569 36159
rect 22569 36125 22603 36159
rect 22603 36125 22612 36159
rect 22560 36116 22612 36125
rect 23756 36252 23808 36304
rect 23480 36184 23532 36236
rect 25320 36184 25372 36236
rect 24400 36159 24452 36168
rect 24400 36125 24409 36159
rect 24409 36125 24443 36159
rect 24443 36125 24452 36159
rect 24400 36116 24452 36125
rect 25504 36116 25556 36168
rect 27436 36320 27488 36372
rect 36544 36320 36596 36372
rect 37096 36252 37148 36304
rect 29460 36184 29512 36236
rect 33784 36227 33836 36236
rect 29000 36116 29052 36168
rect 30012 36116 30064 36168
rect 30196 36159 30248 36168
rect 30196 36125 30205 36159
rect 30205 36125 30239 36159
rect 30239 36125 30248 36159
rect 30196 36116 30248 36125
rect 33784 36193 33793 36227
rect 33793 36193 33827 36227
rect 33827 36193 33836 36227
rect 33784 36184 33836 36193
rect 32404 36116 32456 36168
rect 34244 36116 34296 36168
rect 21272 36048 21324 36100
rect 21732 36091 21784 36100
rect 21732 36057 21741 36091
rect 21741 36057 21775 36091
rect 21775 36057 21784 36091
rect 21732 36048 21784 36057
rect 22100 36048 22152 36100
rect 25964 36048 26016 36100
rect 26240 36091 26292 36100
rect 26240 36057 26258 36091
rect 26258 36057 26292 36091
rect 26240 36048 26292 36057
rect 30288 36048 30340 36100
rect 31852 36048 31904 36100
rect 35440 36091 35492 36100
rect 35440 36057 35474 36091
rect 35474 36057 35492 36091
rect 35440 36048 35492 36057
rect 36084 36048 36136 36100
rect 37740 36159 37792 36168
rect 37740 36125 37749 36159
rect 37749 36125 37783 36159
rect 37783 36125 37792 36159
rect 37740 36116 37792 36125
rect 4712 35980 4764 36032
rect 5080 36023 5132 36032
rect 5080 35989 5089 36023
rect 5089 35989 5123 36023
rect 5123 35989 5132 36023
rect 5080 35980 5132 35989
rect 8208 35980 8260 36032
rect 11428 35980 11480 36032
rect 12072 35980 12124 36032
rect 12624 35980 12676 36032
rect 13268 35980 13320 36032
rect 15844 36023 15896 36032
rect 15844 35989 15853 36023
rect 15853 35989 15887 36023
rect 15887 35989 15896 36023
rect 15844 35980 15896 35989
rect 16304 35980 16356 36032
rect 21088 35980 21140 36032
rect 24584 36023 24636 36032
rect 24584 35989 24593 36023
rect 24593 35989 24627 36023
rect 24627 35989 24636 36023
rect 24584 35980 24636 35989
rect 24860 35980 24912 36032
rect 25228 35980 25280 36032
rect 27712 35980 27764 36032
rect 31668 35980 31720 36032
rect 36544 36023 36596 36032
rect 36544 35989 36553 36023
rect 36553 35989 36587 36023
rect 36587 35989 36596 36023
rect 36544 35980 36596 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 17224 35819 17276 35828
rect 17224 35785 17233 35819
rect 17233 35785 17267 35819
rect 17267 35785 17276 35819
rect 17224 35776 17276 35785
rect 17960 35776 18012 35828
rect 19340 35776 19392 35828
rect 21088 35819 21140 35828
rect 21088 35785 21097 35819
rect 21097 35785 21131 35819
rect 21131 35785 21140 35819
rect 21088 35776 21140 35785
rect 22100 35819 22152 35828
rect 22100 35785 22109 35819
rect 22109 35785 22143 35819
rect 22143 35785 22152 35819
rect 22560 35819 22612 35828
rect 22100 35776 22152 35785
rect 22560 35785 22569 35819
rect 22569 35785 22603 35819
rect 22603 35785 22612 35819
rect 22560 35776 22612 35785
rect 24400 35776 24452 35828
rect 13452 35708 13504 35760
rect 13728 35683 13780 35692
rect 13728 35649 13737 35683
rect 13737 35649 13771 35683
rect 13771 35649 13780 35683
rect 13728 35640 13780 35649
rect 16212 35640 16264 35692
rect 11888 35572 11940 35624
rect 14740 35615 14792 35624
rect 14740 35581 14749 35615
rect 14749 35581 14783 35615
rect 14783 35581 14792 35615
rect 14740 35572 14792 35581
rect 14832 35615 14884 35624
rect 14832 35581 14841 35615
rect 14841 35581 14875 35615
rect 14875 35581 14884 35615
rect 14832 35572 14884 35581
rect 16672 35572 16724 35624
rect 19340 35683 19392 35692
rect 19340 35649 19349 35683
rect 19349 35649 19383 35683
rect 19383 35649 19392 35683
rect 19340 35640 19392 35649
rect 19984 35640 20036 35692
rect 20444 35640 20496 35692
rect 19432 35504 19484 35556
rect 8576 35479 8628 35488
rect 8576 35445 8585 35479
rect 8585 35445 8619 35479
rect 8619 35445 8628 35479
rect 8576 35436 8628 35445
rect 11060 35436 11112 35488
rect 13544 35479 13596 35488
rect 13544 35445 13553 35479
rect 13553 35445 13587 35479
rect 13587 35445 13596 35479
rect 13544 35436 13596 35445
rect 14004 35436 14056 35488
rect 16488 35436 16540 35488
rect 19800 35436 19852 35488
rect 21088 35436 21140 35488
rect 22744 35640 22796 35692
rect 21548 35572 21600 35624
rect 23112 35615 23164 35624
rect 23112 35581 23121 35615
rect 23121 35581 23155 35615
rect 23155 35581 23164 35615
rect 23112 35572 23164 35581
rect 25044 35708 25096 35760
rect 23388 35683 23440 35692
rect 23388 35649 23397 35683
rect 23397 35649 23431 35683
rect 23431 35649 23440 35683
rect 23388 35640 23440 35649
rect 30380 35776 30432 35828
rect 26056 35708 26108 35760
rect 25320 35683 25372 35692
rect 25320 35649 25338 35683
rect 25338 35649 25372 35683
rect 25320 35640 25372 35649
rect 25504 35640 25556 35692
rect 25688 35640 25740 35692
rect 27896 35640 27948 35692
rect 27988 35640 28040 35692
rect 30012 35572 30064 35624
rect 32680 35776 32732 35828
rect 33232 35776 33284 35828
rect 33876 35776 33928 35828
rect 35992 35776 36044 35828
rect 37648 35776 37700 35828
rect 34060 35572 34112 35624
rect 36176 35640 36228 35692
rect 35348 35572 35400 35624
rect 36728 35640 36780 35692
rect 37648 35640 37700 35692
rect 32864 35504 32916 35556
rect 24860 35436 24912 35488
rect 26056 35479 26108 35488
rect 26056 35445 26065 35479
rect 26065 35445 26099 35479
rect 26099 35445 26108 35479
rect 26056 35436 26108 35445
rect 27620 35436 27672 35488
rect 30104 35479 30156 35488
rect 30104 35445 30113 35479
rect 30113 35445 30147 35479
rect 30147 35445 30156 35479
rect 30104 35436 30156 35445
rect 31116 35479 31168 35488
rect 31116 35445 31125 35479
rect 31125 35445 31159 35479
rect 31159 35445 31168 35479
rect 31116 35436 31168 35445
rect 32128 35479 32180 35488
rect 32128 35445 32137 35479
rect 32137 35445 32171 35479
rect 32171 35445 32180 35479
rect 32128 35436 32180 35445
rect 34704 35436 34756 35488
rect 35900 35436 35952 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 10876 35232 10928 35284
rect 13820 35164 13872 35216
rect 14740 35232 14792 35284
rect 19340 35275 19392 35284
rect 15660 35164 15712 35216
rect 12900 35096 12952 35148
rect 16212 35164 16264 35216
rect 6828 35028 6880 35080
rect 14004 35028 14056 35080
rect 14832 35028 14884 35080
rect 15660 35028 15712 35080
rect 19340 35241 19349 35275
rect 19349 35241 19383 35275
rect 19383 35241 19392 35275
rect 19340 35232 19392 35241
rect 23664 35232 23716 35284
rect 25320 35232 25372 35284
rect 26148 35232 26200 35284
rect 27896 35275 27948 35284
rect 27896 35241 27905 35275
rect 27905 35241 27939 35275
rect 27939 35241 27948 35275
rect 27896 35232 27948 35241
rect 16488 35164 16540 35216
rect 16672 35164 16724 35216
rect 20628 35164 20680 35216
rect 22744 35207 22796 35216
rect 22744 35173 22753 35207
rect 22753 35173 22787 35207
rect 22787 35173 22796 35207
rect 22744 35164 22796 35173
rect 23020 35164 23072 35216
rect 25228 35164 25280 35216
rect 25412 35164 25464 35216
rect 27712 35164 27764 35216
rect 31392 35207 31444 35216
rect 31392 35173 31401 35207
rect 31401 35173 31435 35207
rect 31435 35173 31444 35207
rect 31392 35164 31444 35173
rect 16396 35139 16448 35148
rect 16396 35105 16405 35139
rect 16405 35105 16439 35139
rect 16439 35105 16448 35139
rect 16396 35096 16448 35105
rect 10140 34960 10192 35012
rect 12440 34960 12492 35012
rect 16764 35028 16816 35080
rect 29092 35096 29144 35148
rect 19800 35071 19852 35080
rect 19800 35037 19809 35071
rect 19809 35037 19843 35071
rect 19843 35037 19852 35071
rect 19800 35028 19852 35037
rect 20628 35028 20680 35080
rect 21272 35028 21324 35080
rect 24492 35028 24544 35080
rect 24952 35028 25004 35080
rect 26608 35028 26660 35080
rect 30012 35071 30064 35080
rect 30012 35037 30021 35071
rect 30021 35037 30055 35071
rect 30055 35037 30064 35071
rect 30012 35028 30064 35037
rect 33508 35071 33560 35080
rect 33508 35037 33517 35071
rect 33517 35037 33551 35071
rect 33551 35037 33560 35071
rect 33508 35028 33560 35037
rect 33784 35028 33836 35080
rect 34060 35071 34112 35080
rect 34060 35037 34069 35071
rect 34069 35037 34103 35071
rect 34103 35037 34112 35071
rect 36084 35071 36136 35080
rect 34060 35028 34112 35037
rect 9680 34892 9732 34944
rect 11704 34892 11756 34944
rect 12164 34892 12216 34944
rect 14648 34935 14700 34944
rect 14648 34901 14657 34935
rect 14657 34901 14691 34935
rect 14691 34901 14700 34935
rect 14648 34892 14700 34901
rect 14740 34892 14792 34944
rect 22008 34960 22060 35012
rect 31944 34960 31996 35012
rect 34520 34960 34572 35012
rect 19984 34935 20036 34944
rect 19984 34901 19993 34935
rect 19993 34901 20027 34935
rect 20027 34901 20036 34935
rect 19984 34892 20036 34901
rect 20720 34892 20772 34944
rect 21640 34892 21692 34944
rect 22284 34892 22336 34944
rect 23388 34892 23440 34944
rect 24492 34935 24544 34944
rect 24492 34901 24501 34935
rect 24501 34901 24535 34935
rect 24535 34901 24544 34935
rect 24492 34892 24544 34901
rect 25136 34935 25188 34944
rect 25136 34901 25145 34935
rect 25145 34901 25179 34935
rect 25179 34901 25188 34935
rect 25136 34892 25188 34901
rect 28172 34892 28224 34944
rect 31300 34892 31352 34944
rect 34612 34892 34664 34944
rect 36084 35037 36093 35071
rect 36093 35037 36127 35071
rect 36127 35037 36136 35071
rect 36084 35028 36136 35037
rect 37832 34960 37884 35012
rect 36728 34892 36780 34944
rect 37648 34892 37700 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 9404 34688 9456 34740
rect 10876 34731 10928 34740
rect 10876 34697 10885 34731
rect 10885 34697 10919 34731
rect 10919 34697 10928 34731
rect 10876 34688 10928 34697
rect 13544 34688 13596 34740
rect 13728 34688 13780 34740
rect 9956 34620 10008 34672
rect 11888 34620 11940 34672
rect 10232 34595 10284 34604
rect 10232 34561 10241 34595
rect 10241 34561 10275 34595
rect 10275 34561 10284 34595
rect 10232 34552 10284 34561
rect 10324 34595 10376 34604
rect 10324 34561 10333 34595
rect 10333 34561 10367 34595
rect 10367 34561 10376 34595
rect 10324 34552 10376 34561
rect 12164 34595 12216 34604
rect 10140 34484 10192 34536
rect 12164 34561 12173 34595
rect 12173 34561 12207 34595
rect 12207 34561 12216 34595
rect 12164 34552 12216 34561
rect 12348 34552 12400 34604
rect 12900 34595 12952 34604
rect 12900 34561 12909 34595
rect 12909 34561 12943 34595
rect 12943 34561 12952 34595
rect 12900 34552 12952 34561
rect 12808 34484 12860 34536
rect 14096 34484 14148 34536
rect 14648 34688 14700 34740
rect 15016 34688 15068 34740
rect 14740 34663 14792 34672
rect 14740 34629 14749 34663
rect 14749 34629 14783 34663
rect 14783 34629 14792 34663
rect 14740 34620 14792 34629
rect 15660 34663 15712 34672
rect 15660 34629 15669 34663
rect 15669 34629 15703 34663
rect 15703 34629 15712 34663
rect 15660 34620 15712 34629
rect 22008 34731 22060 34740
rect 20444 34620 20496 34672
rect 14924 34595 14976 34604
rect 14924 34561 14933 34595
rect 14933 34561 14967 34595
rect 14967 34561 14976 34595
rect 14924 34552 14976 34561
rect 20720 34620 20772 34672
rect 15200 34484 15252 34536
rect 19432 34484 19484 34536
rect 20260 34484 20312 34536
rect 22008 34697 22017 34731
rect 22017 34697 22051 34731
rect 22051 34697 22060 34731
rect 22008 34688 22060 34697
rect 23388 34731 23440 34740
rect 23388 34697 23397 34731
rect 23397 34697 23431 34731
rect 23431 34697 23440 34731
rect 23388 34688 23440 34697
rect 24308 34731 24360 34740
rect 24308 34697 24317 34731
rect 24317 34697 24351 34731
rect 24351 34697 24360 34731
rect 24308 34688 24360 34697
rect 26240 34731 26292 34740
rect 26240 34697 26249 34731
rect 26249 34697 26283 34731
rect 26283 34697 26292 34731
rect 26240 34688 26292 34697
rect 26976 34731 27028 34740
rect 26976 34697 26985 34731
rect 26985 34697 27019 34731
rect 27019 34697 27028 34731
rect 26976 34688 27028 34697
rect 29092 34731 29144 34740
rect 29092 34697 29101 34731
rect 29101 34697 29135 34731
rect 29135 34697 29144 34731
rect 29092 34688 29144 34697
rect 29184 34688 29236 34740
rect 27988 34620 28040 34672
rect 29644 34620 29696 34672
rect 30012 34620 30064 34672
rect 22560 34595 22612 34604
rect 22560 34561 22569 34595
rect 22569 34561 22603 34595
rect 22603 34561 22612 34595
rect 22560 34552 22612 34561
rect 23204 34595 23256 34604
rect 23204 34561 23213 34595
rect 23213 34561 23247 34595
rect 23247 34561 23256 34595
rect 23204 34552 23256 34561
rect 24860 34552 24912 34604
rect 25596 34552 25648 34604
rect 28080 34595 28132 34604
rect 28080 34561 28098 34595
rect 28098 34561 28132 34595
rect 28080 34552 28132 34561
rect 30196 34595 30248 34604
rect 30196 34561 30214 34595
rect 30214 34561 30248 34595
rect 30196 34552 30248 34561
rect 34796 34552 34848 34604
rect 38200 34552 38252 34604
rect 13084 34416 13136 34468
rect 14924 34416 14976 34468
rect 21640 34484 21692 34536
rect 20904 34416 20956 34468
rect 12992 34391 13044 34400
rect 12992 34357 13001 34391
rect 13001 34357 13035 34391
rect 13035 34357 13044 34391
rect 12992 34348 13044 34357
rect 16580 34348 16632 34400
rect 16856 34348 16908 34400
rect 33048 34391 33100 34400
rect 33048 34357 33057 34391
rect 33057 34357 33091 34391
rect 33091 34357 33100 34391
rect 33048 34348 33100 34357
rect 33140 34348 33192 34400
rect 33508 34348 33560 34400
rect 35992 34484 36044 34536
rect 36268 34459 36320 34468
rect 36268 34425 36277 34459
rect 36277 34425 36311 34459
rect 36311 34425 36320 34459
rect 36268 34416 36320 34425
rect 36360 34391 36412 34400
rect 36360 34357 36369 34391
rect 36369 34357 36403 34391
rect 36403 34357 36412 34391
rect 36360 34348 36412 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 10324 34144 10376 34196
rect 12256 34119 12308 34128
rect 12256 34085 12265 34119
rect 12265 34085 12299 34119
rect 12299 34085 12308 34119
rect 12256 34076 12308 34085
rect 15108 34144 15160 34196
rect 16672 34187 16724 34196
rect 16672 34153 16681 34187
rect 16681 34153 16715 34187
rect 16715 34153 16724 34187
rect 22192 34187 22244 34196
rect 16672 34144 16724 34153
rect 22192 34153 22201 34187
rect 22201 34153 22235 34187
rect 22235 34153 22244 34187
rect 22192 34144 22244 34153
rect 23204 34144 23256 34196
rect 24952 34187 25004 34196
rect 24952 34153 24961 34187
rect 24961 34153 24995 34187
rect 24995 34153 25004 34187
rect 24952 34144 25004 34153
rect 25412 34144 25464 34196
rect 25780 34144 25832 34196
rect 29000 34187 29052 34196
rect 29000 34153 29009 34187
rect 29009 34153 29043 34187
rect 29043 34153 29052 34187
rect 29000 34144 29052 34153
rect 30196 34144 30248 34196
rect 16396 34076 16448 34128
rect 12992 34008 13044 34060
rect 14924 34008 14976 34060
rect 9220 33983 9272 33992
rect 9220 33949 9229 33983
rect 9229 33949 9263 33983
rect 9263 33949 9272 33983
rect 9220 33940 9272 33949
rect 9404 33983 9456 33992
rect 9404 33949 9413 33983
rect 9413 33949 9447 33983
rect 9447 33949 9456 33983
rect 9404 33940 9456 33949
rect 10232 33940 10284 33992
rect 11888 33940 11940 33992
rect 13820 33940 13872 33992
rect 14096 33983 14148 33992
rect 14096 33949 14105 33983
rect 14105 33949 14139 33983
rect 14139 33949 14148 33983
rect 14096 33940 14148 33949
rect 17684 33983 17736 33992
rect 12900 33872 12952 33924
rect 17684 33949 17693 33983
rect 17693 33949 17727 33983
rect 17727 33949 17736 33983
rect 17684 33940 17736 33949
rect 22100 34008 22152 34060
rect 23204 34008 23256 34060
rect 24584 34008 24636 34060
rect 24768 34008 24820 34060
rect 29644 34008 29696 34060
rect 15016 33915 15068 33924
rect 15016 33881 15025 33915
rect 15025 33881 15059 33915
rect 15059 33881 15068 33915
rect 15016 33872 15068 33881
rect 15200 33915 15252 33924
rect 15200 33881 15225 33915
rect 15225 33881 15252 33915
rect 15200 33872 15252 33881
rect 16488 33872 16540 33924
rect 16580 33915 16632 33924
rect 16580 33881 16589 33915
rect 16589 33881 16623 33915
rect 16623 33881 16632 33915
rect 16580 33872 16632 33881
rect 16672 33804 16724 33856
rect 18328 33915 18380 33924
rect 18328 33881 18337 33915
rect 18337 33881 18371 33915
rect 18371 33881 18380 33915
rect 18328 33872 18380 33881
rect 20444 33940 20496 33992
rect 21824 33940 21876 33992
rect 25136 33940 25188 33992
rect 27804 33983 27856 33992
rect 27804 33949 27822 33983
rect 27822 33949 27856 33983
rect 27804 33940 27856 33949
rect 35992 34144 36044 34196
rect 35900 33940 35952 33992
rect 36084 33940 36136 33992
rect 33232 33872 33284 33924
rect 34520 33872 34572 33924
rect 18052 33804 18104 33856
rect 23112 33804 23164 33856
rect 24032 33804 24084 33856
rect 24584 33804 24636 33856
rect 33140 33804 33192 33856
rect 34244 33804 34296 33856
rect 37096 33872 37148 33924
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 8760 33643 8812 33652
rect 8760 33609 8769 33643
rect 8769 33609 8803 33643
rect 8803 33609 8812 33643
rect 8760 33600 8812 33609
rect 10232 33600 10284 33652
rect 13084 33600 13136 33652
rect 13176 33600 13228 33652
rect 13360 33600 13412 33652
rect 20076 33600 20128 33652
rect 20444 33643 20496 33652
rect 20444 33609 20453 33643
rect 20453 33609 20487 33643
rect 20487 33609 20496 33643
rect 20444 33600 20496 33609
rect 21824 33643 21876 33652
rect 21824 33609 21833 33643
rect 21833 33609 21867 33643
rect 21867 33609 21876 33643
rect 21824 33600 21876 33609
rect 22560 33600 22612 33652
rect 24492 33600 24544 33652
rect 37740 33600 37792 33652
rect 8852 33464 8904 33516
rect 9680 33464 9732 33516
rect 9220 33396 9272 33448
rect 13820 33532 13872 33584
rect 26056 33532 26108 33584
rect 12808 33507 12860 33516
rect 12808 33473 12817 33507
rect 12817 33473 12851 33507
rect 12851 33473 12860 33507
rect 12808 33464 12860 33473
rect 13176 33464 13228 33516
rect 14096 33464 14148 33516
rect 16672 33507 16724 33516
rect 16672 33473 16681 33507
rect 16681 33473 16715 33507
rect 16715 33473 16724 33507
rect 16672 33464 16724 33473
rect 18236 33507 18288 33516
rect 18236 33473 18245 33507
rect 18245 33473 18279 33507
rect 18279 33473 18288 33507
rect 18236 33464 18288 33473
rect 20076 33507 20128 33516
rect 20076 33473 20085 33507
rect 20085 33473 20119 33507
rect 20119 33473 20128 33507
rect 20076 33464 20128 33473
rect 22744 33464 22796 33516
rect 22928 33464 22980 33516
rect 27620 33464 27672 33516
rect 27804 33464 27856 33516
rect 33232 33464 33284 33516
rect 36360 33464 36412 33516
rect 18052 33396 18104 33448
rect 20628 33396 20680 33448
rect 23204 33396 23256 33448
rect 35900 33396 35952 33448
rect 23664 33328 23716 33380
rect 12716 33260 12768 33312
rect 14372 33260 14424 33312
rect 15108 33260 15160 33312
rect 16764 33260 16816 33312
rect 17684 33260 17736 33312
rect 18144 33260 18196 33312
rect 20812 33260 20864 33312
rect 29644 33260 29696 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 9680 33056 9732 33108
rect 12348 33056 12400 33108
rect 18236 33056 18288 33108
rect 22100 33056 22152 33108
rect 18052 32988 18104 33040
rect 22744 33031 22796 33040
rect 22744 32997 22753 33031
rect 22753 32997 22787 33031
rect 22787 32997 22796 33031
rect 22744 32988 22796 32997
rect 23296 33031 23348 33040
rect 23296 32997 23305 33031
rect 23305 32997 23339 33031
rect 23339 32997 23348 33031
rect 23296 32988 23348 32997
rect 24400 33031 24452 33040
rect 24400 32997 24409 33031
rect 24409 32997 24443 33031
rect 24443 32997 24452 33031
rect 24400 32988 24452 32997
rect 17868 32920 17920 32972
rect 20076 32920 20128 32972
rect 22100 32920 22152 32972
rect 12716 32852 12768 32904
rect 12900 32852 12952 32904
rect 19248 32852 19300 32904
rect 19156 32784 19208 32836
rect 25780 32895 25832 32904
rect 25780 32861 25789 32895
rect 25789 32861 25823 32895
rect 25823 32861 25832 32895
rect 25780 32852 25832 32861
rect 26056 32852 26108 32904
rect 29000 32852 29052 32904
rect 33140 32852 33192 32904
rect 21364 32784 21416 32836
rect 24400 32784 24452 32836
rect 24492 32784 24544 32836
rect 14188 32759 14240 32768
rect 14188 32725 14197 32759
rect 14197 32725 14231 32759
rect 14231 32725 14240 32759
rect 14188 32716 14240 32725
rect 23112 32716 23164 32768
rect 27252 32784 27304 32836
rect 33324 32784 33376 32836
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 5080 32444 5132 32496
rect 12900 32444 12952 32496
rect 13176 32487 13228 32496
rect 13176 32453 13185 32487
rect 13185 32453 13219 32487
rect 13219 32453 13228 32487
rect 13176 32444 13228 32453
rect 12256 32419 12308 32428
rect 12256 32385 12265 32419
rect 12265 32385 12299 32419
rect 12299 32385 12308 32419
rect 12256 32376 12308 32385
rect 14188 32444 14240 32496
rect 13912 32419 13964 32428
rect 13912 32385 13921 32419
rect 13921 32385 13955 32419
rect 13955 32385 13964 32419
rect 13912 32376 13964 32385
rect 15016 32444 15068 32496
rect 23388 32444 23440 32496
rect 36268 32512 36320 32564
rect 16764 32376 16816 32428
rect 22468 32376 22520 32428
rect 26056 32419 26108 32428
rect 18788 32351 18840 32360
rect 18788 32317 18797 32351
rect 18797 32317 18831 32351
rect 18831 32317 18840 32351
rect 18788 32308 18840 32317
rect 16580 32240 16632 32292
rect 17040 32240 17092 32292
rect 22744 32240 22796 32292
rect 26056 32385 26065 32419
rect 26065 32385 26099 32419
rect 26099 32385 26108 32419
rect 26056 32376 26108 32385
rect 26148 32376 26200 32428
rect 29736 32376 29788 32428
rect 29644 32351 29696 32360
rect 29644 32317 29653 32351
rect 29653 32317 29687 32351
rect 29687 32317 29696 32351
rect 29644 32308 29696 32317
rect 31024 32283 31076 32292
rect 31024 32249 31033 32283
rect 31033 32249 31067 32283
rect 31067 32249 31076 32283
rect 31024 32240 31076 32249
rect 13912 32172 13964 32224
rect 15936 32172 15988 32224
rect 16488 32172 16540 32224
rect 21456 32172 21508 32224
rect 24676 32215 24728 32224
rect 24676 32181 24685 32215
rect 24685 32181 24719 32215
rect 24719 32181 24728 32215
rect 24676 32172 24728 32181
rect 27620 32172 27672 32224
rect 35900 32172 35952 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 13912 31968 13964 32020
rect 15016 31968 15068 32020
rect 21364 31900 21416 31952
rect 26148 31968 26200 32020
rect 29552 31968 29604 32020
rect 29736 31968 29788 32020
rect 31392 31968 31444 32020
rect 34796 32011 34848 32020
rect 24400 31943 24452 31952
rect 15936 31875 15988 31884
rect 15936 31841 15945 31875
rect 15945 31841 15979 31875
rect 15979 31841 15988 31875
rect 15936 31832 15988 31841
rect 17132 31832 17184 31884
rect 20720 31832 20772 31884
rect 21088 31875 21140 31884
rect 21088 31841 21097 31875
rect 21097 31841 21131 31875
rect 21131 31841 21140 31875
rect 21088 31832 21140 31841
rect 24400 31909 24409 31943
rect 24409 31909 24443 31943
rect 24443 31909 24452 31943
rect 24400 31900 24452 31909
rect 31208 31900 31260 31952
rect 16304 31764 16356 31816
rect 18788 31764 18840 31816
rect 22008 31807 22060 31816
rect 21456 31696 21508 31748
rect 22008 31773 22017 31807
rect 22017 31773 22051 31807
rect 22051 31773 22060 31807
rect 22008 31764 22060 31773
rect 24768 31832 24820 31884
rect 26056 31832 26108 31884
rect 24952 31764 25004 31816
rect 25044 31764 25096 31816
rect 33140 31764 33192 31816
rect 34796 31977 34805 32011
rect 34805 31977 34839 32011
rect 34839 31977 34848 32011
rect 34796 31968 34848 31977
rect 34704 31900 34756 31952
rect 35900 31832 35952 31884
rect 23112 31671 23164 31680
rect 23112 31637 23121 31671
rect 23121 31637 23155 31671
rect 23155 31637 23164 31671
rect 23112 31628 23164 31637
rect 30656 31628 30708 31680
rect 35256 31671 35308 31680
rect 35256 31637 35265 31671
rect 35265 31637 35299 31671
rect 35299 31637 35308 31671
rect 35256 31628 35308 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 16672 31331 16724 31340
rect 16672 31297 16681 31331
rect 16681 31297 16715 31331
rect 16715 31297 16724 31331
rect 16672 31288 16724 31297
rect 27620 31424 27672 31476
rect 34888 31424 34940 31476
rect 35624 31424 35676 31476
rect 20352 31356 20404 31408
rect 23112 31356 23164 31408
rect 25596 31356 25648 31408
rect 29644 31356 29696 31408
rect 20444 31331 20496 31340
rect 20444 31297 20453 31331
rect 20453 31297 20487 31331
rect 20487 31297 20496 31331
rect 20444 31288 20496 31297
rect 24400 31288 24452 31340
rect 26056 31288 26108 31340
rect 29000 31288 29052 31340
rect 34796 31356 34848 31408
rect 33140 31288 33192 31340
rect 17040 31220 17092 31272
rect 20720 31220 20772 31272
rect 20812 31220 20864 31272
rect 21916 31263 21968 31272
rect 21916 31229 21925 31263
rect 21925 31229 21959 31263
rect 21959 31229 21968 31263
rect 21916 31220 21968 31229
rect 4712 31152 4764 31204
rect 17776 31084 17828 31136
rect 17960 31127 18012 31136
rect 17960 31093 17969 31127
rect 17969 31093 18003 31127
rect 18003 31093 18012 31127
rect 17960 31084 18012 31093
rect 18144 31084 18196 31136
rect 24492 31152 24544 31204
rect 34612 31220 34664 31272
rect 35256 31288 35308 31340
rect 22560 31127 22612 31136
rect 22560 31093 22569 31127
rect 22569 31093 22603 31127
rect 22603 31093 22612 31127
rect 22560 31084 22612 31093
rect 24308 31127 24360 31136
rect 24308 31093 24317 31127
rect 24317 31093 24351 31127
rect 24351 31093 24360 31127
rect 24308 31084 24360 31093
rect 28080 31084 28132 31136
rect 28356 31127 28408 31136
rect 28356 31093 28365 31127
rect 28365 31093 28399 31127
rect 28399 31093 28408 31127
rect 28356 31084 28408 31093
rect 29092 31127 29144 31136
rect 29092 31093 29101 31127
rect 29101 31093 29135 31127
rect 29135 31093 29144 31127
rect 29092 31084 29144 31093
rect 33140 31084 33192 31136
rect 36084 31127 36136 31136
rect 36084 31093 36093 31127
rect 36093 31093 36127 31127
rect 36127 31093 36136 31127
rect 36084 31084 36136 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 12256 30880 12308 30932
rect 17776 30880 17828 30932
rect 18052 30812 18104 30864
rect 20444 30880 20496 30932
rect 22008 30880 22060 30932
rect 32128 30880 32180 30932
rect 36452 30923 36504 30932
rect 36452 30889 36461 30923
rect 36461 30889 36495 30923
rect 36495 30889 36504 30923
rect 36452 30880 36504 30889
rect 19984 30812 20036 30864
rect 21548 30812 21600 30864
rect 24308 30812 24360 30864
rect 17132 30787 17184 30796
rect 17132 30753 17141 30787
rect 17141 30753 17175 30787
rect 17175 30753 17184 30787
rect 26056 30787 26108 30796
rect 17132 30744 17184 30753
rect 11796 30719 11848 30728
rect 11796 30685 11805 30719
rect 11805 30685 11839 30719
rect 11839 30685 11848 30719
rect 11796 30676 11848 30685
rect 11980 30719 12032 30728
rect 11980 30685 11989 30719
rect 11989 30685 12023 30719
rect 12023 30685 12032 30719
rect 11980 30676 12032 30685
rect 12624 30719 12676 30728
rect 12624 30685 12633 30719
rect 12633 30685 12667 30719
rect 12667 30685 12676 30719
rect 12624 30676 12676 30685
rect 17960 30676 18012 30728
rect 26056 30753 26065 30787
rect 26065 30753 26099 30787
rect 26099 30753 26108 30787
rect 26056 30744 26108 30753
rect 20536 30719 20588 30728
rect 18052 30608 18104 30660
rect 20536 30685 20545 30719
rect 20545 30685 20579 30719
rect 20579 30685 20588 30719
rect 20536 30676 20588 30685
rect 20720 30719 20772 30728
rect 20720 30685 20729 30719
rect 20729 30685 20763 30719
rect 20763 30685 20772 30719
rect 20720 30676 20772 30685
rect 27804 30719 27856 30728
rect 27804 30685 27813 30719
rect 27813 30685 27847 30719
rect 27847 30685 27856 30719
rect 27804 30676 27856 30685
rect 32312 30719 32364 30728
rect 32312 30685 32321 30719
rect 32321 30685 32355 30719
rect 32355 30685 32364 30719
rect 32312 30676 32364 30685
rect 35900 30676 35952 30728
rect 12808 30583 12860 30592
rect 12808 30549 12817 30583
rect 12817 30549 12851 30583
rect 12851 30549 12860 30583
rect 12808 30540 12860 30549
rect 17592 30583 17644 30592
rect 17592 30549 17601 30583
rect 17601 30549 17635 30583
rect 17635 30549 17644 30583
rect 17592 30540 17644 30549
rect 35716 30608 35768 30660
rect 32128 30540 32180 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 12808 30336 12860 30388
rect 12624 30268 12676 30320
rect 16672 30268 16724 30320
rect 20536 30268 20588 30320
rect 22192 30268 22244 30320
rect 12256 30200 12308 30252
rect 14372 30243 14424 30252
rect 14372 30209 14381 30243
rect 14381 30209 14415 30243
rect 14415 30209 14424 30243
rect 14372 30200 14424 30209
rect 15016 30200 15068 30252
rect 15292 30243 15344 30252
rect 15292 30209 15301 30243
rect 15301 30209 15335 30243
rect 15335 30209 15344 30243
rect 15292 30200 15344 30209
rect 17500 30243 17552 30252
rect 17500 30209 17509 30243
rect 17509 30209 17543 30243
rect 17543 30209 17552 30243
rect 17500 30200 17552 30209
rect 21732 30200 21784 30252
rect 29000 30268 29052 30320
rect 27620 30200 27672 30252
rect 28356 30200 28408 30252
rect 33416 30200 33468 30252
rect 11796 30132 11848 30184
rect 12624 29996 12676 30048
rect 15200 30132 15252 30184
rect 26516 30132 26568 30184
rect 14372 29996 14424 30048
rect 18052 29996 18104 30048
rect 18604 29996 18656 30048
rect 22100 29996 22152 30048
rect 24400 30039 24452 30048
rect 24400 30005 24409 30039
rect 24409 30005 24443 30039
rect 24443 30005 24452 30039
rect 24400 29996 24452 30005
rect 25872 30064 25924 30116
rect 26332 30064 26384 30116
rect 25596 29996 25648 30048
rect 26424 29996 26476 30048
rect 35900 30132 35952 30184
rect 29276 29996 29328 30048
rect 30288 30039 30340 30048
rect 30288 30005 30297 30039
rect 30297 30005 30331 30039
rect 30331 30005 30340 30039
rect 30288 29996 30340 30005
rect 33508 30039 33560 30048
rect 33508 30005 33517 30039
rect 33517 30005 33551 30039
rect 33551 30005 33560 30039
rect 33508 29996 33560 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 11980 29792 12032 29844
rect 16488 29835 16540 29844
rect 16488 29801 16497 29835
rect 16497 29801 16531 29835
rect 16531 29801 16540 29835
rect 16488 29792 16540 29801
rect 13544 29767 13596 29776
rect 13544 29733 13553 29767
rect 13553 29733 13587 29767
rect 13587 29733 13596 29767
rect 13544 29724 13596 29733
rect 13728 29724 13780 29776
rect 24400 29792 24452 29844
rect 25136 29792 25188 29844
rect 25964 29792 26016 29844
rect 30288 29792 30340 29844
rect 22008 29767 22060 29776
rect 12808 29699 12860 29708
rect 12808 29665 12817 29699
rect 12817 29665 12851 29699
rect 12851 29665 12860 29699
rect 12808 29656 12860 29665
rect 15936 29656 15988 29708
rect 22008 29733 22017 29767
rect 22017 29733 22051 29767
rect 22051 29733 22060 29767
rect 22008 29724 22060 29733
rect 28908 29724 28960 29776
rect 33508 29792 33560 29844
rect 36176 29792 36228 29844
rect 37924 29792 37976 29844
rect 38108 29835 38160 29844
rect 38108 29801 38117 29835
rect 38117 29801 38151 29835
rect 38151 29801 38160 29835
rect 38108 29792 38160 29801
rect 21732 29656 21784 29708
rect 22192 29656 22244 29708
rect 12624 29588 12676 29640
rect 14096 29631 14148 29640
rect 14096 29597 14105 29631
rect 14105 29597 14139 29631
rect 14139 29597 14148 29631
rect 14096 29588 14148 29597
rect 16488 29588 16540 29640
rect 17592 29588 17644 29640
rect 21088 29631 21140 29640
rect 21088 29597 21097 29631
rect 21097 29597 21131 29631
rect 21131 29597 21140 29631
rect 21088 29588 21140 29597
rect 22100 29631 22152 29640
rect 22100 29597 22108 29631
rect 22108 29597 22142 29631
rect 22142 29597 22152 29631
rect 22560 29631 22612 29640
rect 22100 29588 22152 29597
rect 22560 29597 22569 29631
rect 22569 29597 22603 29631
rect 22603 29597 22612 29631
rect 22560 29588 22612 29597
rect 32312 29656 32364 29708
rect 10140 29520 10192 29572
rect 20996 29520 21048 29572
rect 24860 29520 24912 29572
rect 26516 29588 26568 29640
rect 35900 29588 35952 29640
rect 29092 29520 29144 29572
rect 12900 29452 12952 29504
rect 13544 29452 13596 29504
rect 14280 29495 14332 29504
rect 14280 29461 14289 29495
rect 14289 29461 14323 29495
rect 14323 29461 14332 29495
rect 14280 29452 14332 29461
rect 15384 29452 15436 29504
rect 15752 29452 15804 29504
rect 17224 29495 17276 29504
rect 17224 29461 17233 29495
rect 17233 29461 17267 29495
rect 17267 29461 17276 29495
rect 17224 29452 17276 29461
rect 22100 29452 22152 29504
rect 22744 29495 22796 29504
rect 22744 29461 22753 29495
rect 22753 29461 22787 29495
rect 22787 29461 22796 29495
rect 22744 29452 22796 29461
rect 24400 29495 24452 29504
rect 24400 29461 24409 29495
rect 24409 29461 24443 29495
rect 24443 29461 24452 29495
rect 24400 29452 24452 29461
rect 28172 29452 28224 29504
rect 35440 29520 35492 29572
rect 36544 29520 36596 29572
rect 31852 29452 31904 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 10140 29248 10192 29300
rect 13176 29291 13228 29300
rect 13176 29257 13185 29291
rect 13185 29257 13219 29291
rect 13219 29257 13228 29291
rect 13176 29248 13228 29257
rect 16304 29248 16356 29300
rect 17224 29248 17276 29300
rect 20812 29223 20864 29232
rect 20812 29189 20821 29223
rect 20821 29189 20855 29223
rect 20855 29189 20864 29223
rect 20812 29180 20864 29189
rect 20996 29180 21048 29232
rect 25596 29248 25648 29300
rect 22744 29180 22796 29232
rect 32312 29180 32364 29232
rect 12164 29155 12216 29164
rect 12164 29121 12173 29155
rect 12173 29121 12207 29155
rect 12207 29121 12216 29155
rect 12164 29112 12216 29121
rect 12992 29155 13044 29164
rect 12992 29121 13001 29155
rect 13001 29121 13035 29155
rect 13035 29121 13044 29155
rect 12992 29112 13044 29121
rect 15384 29155 15436 29164
rect 15384 29121 15393 29155
rect 15393 29121 15427 29155
rect 15427 29121 15436 29155
rect 15384 29112 15436 29121
rect 19340 29112 19392 29164
rect 21824 29155 21876 29164
rect 21824 29121 21833 29155
rect 21833 29121 21867 29155
rect 21867 29121 21876 29155
rect 21824 29112 21876 29121
rect 22008 29155 22060 29164
rect 22008 29121 22017 29155
rect 22017 29121 22051 29155
rect 22051 29121 22060 29155
rect 22008 29112 22060 29121
rect 22468 29112 22520 29164
rect 8576 29044 8628 29096
rect 12532 29044 12584 29096
rect 13728 29044 13780 29096
rect 15200 29087 15252 29096
rect 15200 29053 15209 29087
rect 15209 29053 15243 29087
rect 15243 29053 15252 29087
rect 15200 29044 15252 29053
rect 21088 29044 21140 29096
rect 10508 28976 10560 29028
rect 12348 29019 12400 29028
rect 12348 28985 12357 29019
rect 12357 28985 12391 29019
rect 12391 28985 12400 29019
rect 12348 28976 12400 28985
rect 15752 28976 15804 29028
rect 29276 29112 29328 29164
rect 30564 29112 30616 29164
rect 26516 29044 26568 29096
rect 24492 28976 24544 29028
rect 27988 29019 28040 29028
rect 27988 28985 27997 29019
rect 27997 28985 28031 29019
rect 28031 28985 28040 29019
rect 27988 28976 28040 28985
rect 32864 29019 32916 29028
rect 32864 28985 32873 29019
rect 32873 28985 32907 29019
rect 32907 28985 32916 29019
rect 32864 28976 32916 28985
rect 9588 28908 9640 28960
rect 10876 28908 10928 28960
rect 21180 28908 21232 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 14096 28747 14148 28756
rect 14096 28713 14105 28747
rect 14105 28713 14139 28747
rect 14139 28713 14148 28747
rect 14096 28704 14148 28713
rect 17500 28704 17552 28756
rect 21824 28704 21876 28756
rect 12072 28636 12124 28688
rect 15660 28636 15712 28688
rect 18604 28636 18656 28688
rect 9588 28568 9640 28620
rect 5816 28500 5868 28552
rect 9128 28500 9180 28552
rect 10508 28500 10560 28552
rect 10876 28500 10928 28552
rect 11612 28543 11664 28552
rect 11612 28509 11621 28543
rect 11621 28509 11655 28543
rect 11655 28509 11664 28543
rect 11612 28500 11664 28509
rect 12348 28475 12400 28484
rect 12348 28441 12357 28475
rect 12357 28441 12391 28475
rect 12391 28441 12400 28475
rect 12348 28432 12400 28441
rect 9036 28407 9088 28416
rect 9036 28373 9045 28407
rect 9045 28373 9079 28407
rect 9079 28373 9088 28407
rect 9036 28364 9088 28373
rect 10048 28364 10100 28416
rect 10232 28407 10284 28416
rect 10232 28373 10241 28407
rect 10241 28373 10275 28407
rect 10275 28373 10284 28407
rect 10232 28364 10284 28373
rect 11796 28407 11848 28416
rect 11796 28373 11805 28407
rect 11805 28373 11839 28407
rect 11839 28373 11848 28407
rect 11796 28364 11848 28373
rect 14280 28543 14332 28552
rect 14280 28509 14289 28543
rect 14289 28509 14323 28543
rect 14323 28509 14332 28543
rect 14280 28500 14332 28509
rect 15016 28475 15068 28484
rect 15016 28441 15025 28475
rect 15025 28441 15059 28475
rect 15059 28441 15068 28475
rect 15016 28432 15068 28441
rect 15200 28475 15252 28484
rect 15200 28441 15209 28475
rect 15209 28441 15243 28475
rect 15243 28441 15252 28475
rect 15200 28432 15252 28441
rect 13820 28364 13872 28416
rect 20536 28568 20588 28620
rect 21088 28568 21140 28620
rect 21824 28611 21876 28620
rect 21824 28577 21833 28611
rect 21833 28577 21867 28611
rect 21867 28577 21876 28611
rect 21824 28568 21876 28577
rect 38016 28704 38068 28756
rect 17224 28543 17276 28552
rect 17224 28509 17233 28543
rect 17233 28509 17267 28543
rect 17267 28509 17276 28543
rect 17224 28500 17276 28509
rect 21180 28543 21232 28552
rect 21180 28509 21189 28543
rect 21189 28509 21223 28543
rect 21223 28509 21232 28543
rect 21180 28500 21232 28509
rect 29276 28568 29328 28620
rect 32312 28611 32364 28620
rect 32312 28577 32321 28611
rect 32321 28577 32355 28611
rect 32355 28577 32364 28611
rect 32312 28568 32364 28577
rect 18788 28432 18840 28484
rect 18880 28432 18932 28484
rect 26516 28500 26568 28552
rect 36820 28500 36872 28552
rect 16212 28407 16264 28416
rect 16212 28373 16221 28407
rect 16221 28373 16255 28407
rect 16255 28373 16264 28407
rect 16212 28364 16264 28373
rect 25596 28432 25648 28484
rect 31760 28432 31812 28484
rect 36176 28432 36228 28484
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 9956 28203 10008 28212
rect 9956 28169 9965 28203
rect 9965 28169 9999 28203
rect 9999 28169 10008 28203
rect 9956 28160 10008 28169
rect 12164 28160 12216 28212
rect 12992 28160 13044 28212
rect 15292 28160 15344 28212
rect 15660 28160 15712 28212
rect 19340 28160 19392 28212
rect 11796 28092 11848 28144
rect 29276 28092 29328 28144
rect 9036 28067 9088 28076
rect 9036 28033 9045 28067
rect 9045 28033 9079 28067
rect 9079 28033 9088 28067
rect 9036 28024 9088 28033
rect 10232 28024 10284 28076
rect 11888 28067 11940 28076
rect 11888 28033 11897 28067
rect 11897 28033 11931 28067
rect 11931 28033 11940 28067
rect 11888 28024 11940 28033
rect 12072 28067 12124 28076
rect 12072 28033 12081 28067
rect 12081 28033 12115 28067
rect 12115 28033 12124 28067
rect 12072 28024 12124 28033
rect 13268 28024 13320 28076
rect 16212 28024 16264 28076
rect 16672 28067 16724 28076
rect 16672 28033 16681 28067
rect 16681 28033 16715 28067
rect 16715 28033 16724 28067
rect 16672 28024 16724 28033
rect 18972 28067 19024 28076
rect 18972 28033 18981 28067
rect 18981 28033 19015 28067
rect 19015 28033 19024 28067
rect 18972 28024 19024 28033
rect 29736 28067 29788 28076
rect 34520 28092 34572 28144
rect 29736 28033 29754 28067
rect 29754 28033 29788 28067
rect 29736 28024 29788 28033
rect 11060 27956 11112 28008
rect 15200 27956 15252 28008
rect 15936 27999 15988 28008
rect 15936 27965 15945 27999
rect 15945 27965 15979 27999
rect 15979 27965 15988 27999
rect 15936 27956 15988 27965
rect 18788 27999 18840 28008
rect 18788 27965 18797 27999
rect 18797 27965 18831 27999
rect 18831 27965 18840 27999
rect 18788 27956 18840 27965
rect 26240 27956 26292 28008
rect 26516 27956 26568 28008
rect 35900 27956 35952 28008
rect 37004 27956 37056 28008
rect 13452 27888 13504 27940
rect 16856 27931 16908 27940
rect 11704 27820 11756 27872
rect 13544 27863 13596 27872
rect 13544 27829 13553 27863
rect 13553 27829 13587 27863
rect 13587 27829 13596 27863
rect 13544 27820 13596 27829
rect 14924 27863 14976 27872
rect 14924 27829 14933 27863
rect 14933 27829 14967 27863
rect 14967 27829 14976 27863
rect 14924 27820 14976 27829
rect 16856 27897 16865 27931
rect 16865 27897 16899 27931
rect 16899 27897 16908 27931
rect 16856 27888 16908 27897
rect 20536 27820 20588 27872
rect 25044 27820 25096 27872
rect 32036 27820 32088 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 11060 27616 11112 27668
rect 11612 27616 11664 27668
rect 12072 27616 12124 27668
rect 16672 27548 16724 27600
rect 18696 27591 18748 27600
rect 12808 27480 12860 27532
rect 13820 27480 13872 27532
rect 14924 27480 14976 27532
rect 15200 27480 15252 27532
rect 16488 27480 16540 27532
rect 18696 27557 18705 27591
rect 18705 27557 18739 27591
rect 18739 27557 18748 27591
rect 18696 27548 18748 27557
rect 19248 27591 19300 27600
rect 19248 27557 19257 27591
rect 19257 27557 19291 27591
rect 19291 27557 19300 27591
rect 19248 27548 19300 27557
rect 11060 27455 11112 27464
rect 11060 27421 11069 27455
rect 11069 27421 11103 27455
rect 11103 27421 11112 27455
rect 11060 27412 11112 27421
rect 11152 27412 11204 27464
rect 15476 27455 15528 27464
rect 10508 27344 10560 27396
rect 13544 27344 13596 27396
rect 15200 27344 15252 27396
rect 7564 27276 7616 27328
rect 14464 27319 14516 27328
rect 14464 27285 14473 27319
rect 14473 27285 14507 27319
rect 14507 27285 14516 27319
rect 14464 27276 14516 27285
rect 14556 27276 14608 27328
rect 15476 27421 15485 27455
rect 15485 27421 15519 27455
rect 15519 27421 15528 27455
rect 15476 27412 15528 27421
rect 15660 27412 15712 27464
rect 17132 27412 17184 27464
rect 18512 27455 18564 27464
rect 18512 27421 18521 27455
rect 18521 27421 18555 27455
rect 18555 27421 18564 27455
rect 18512 27412 18564 27421
rect 17868 27276 17920 27328
rect 20812 27412 20864 27464
rect 22560 27412 22612 27464
rect 26424 27480 26476 27532
rect 26240 27412 26292 27464
rect 30104 27548 30156 27600
rect 29276 27480 29328 27532
rect 29368 27480 29420 27532
rect 30196 27480 30248 27532
rect 30656 27412 30708 27464
rect 31760 27412 31812 27464
rect 31944 27412 31996 27464
rect 32312 27412 32364 27464
rect 33048 27412 33100 27464
rect 37004 27455 37056 27464
rect 37004 27421 37013 27455
rect 37013 27421 37047 27455
rect 37047 27421 37056 27455
rect 37004 27412 37056 27421
rect 20720 27344 20772 27396
rect 24860 27344 24912 27396
rect 26424 27344 26476 27396
rect 30748 27344 30800 27396
rect 20536 27276 20588 27328
rect 21824 27319 21876 27328
rect 21824 27285 21833 27319
rect 21833 27285 21867 27319
rect 21867 27285 21876 27319
rect 21824 27276 21876 27285
rect 24308 27276 24360 27328
rect 24400 27319 24452 27328
rect 24400 27285 24409 27319
rect 24409 27285 24443 27319
rect 24443 27285 24452 27319
rect 24400 27276 24452 27285
rect 25044 27276 25096 27328
rect 30472 27276 30524 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 12256 27072 12308 27124
rect 12532 27072 12584 27124
rect 18512 27072 18564 27124
rect 20812 27115 20864 27124
rect 20812 27081 20821 27115
rect 20821 27081 20855 27115
rect 20855 27081 20864 27115
rect 20812 27072 20864 27081
rect 21824 27072 21876 27124
rect 31484 27072 31536 27124
rect 35348 27115 35400 27124
rect 35348 27081 35357 27115
rect 35357 27081 35391 27115
rect 35391 27081 35400 27115
rect 35348 27072 35400 27081
rect 35624 27072 35676 27124
rect 14464 27004 14516 27056
rect 8576 26979 8628 26988
rect 8576 26945 8585 26979
rect 8585 26945 8619 26979
rect 8619 26945 8628 26979
rect 8576 26936 8628 26945
rect 9128 26936 9180 26988
rect 11244 26936 11296 26988
rect 13176 26936 13228 26988
rect 14372 26979 14424 26988
rect 14372 26945 14381 26979
rect 14381 26945 14415 26979
rect 14415 26945 14424 26979
rect 14372 26936 14424 26945
rect 14556 26979 14608 26988
rect 14556 26945 14565 26979
rect 14565 26945 14599 26979
rect 14599 26945 14608 26979
rect 14556 26936 14608 26945
rect 14924 26936 14976 26988
rect 16948 26936 17000 26988
rect 17592 26979 17644 26988
rect 17592 26945 17601 26979
rect 17601 26945 17635 26979
rect 17635 26945 17644 26979
rect 17592 26936 17644 26945
rect 17868 27004 17920 27056
rect 22560 27004 22612 27056
rect 22652 27004 22704 27056
rect 31116 27004 31168 27056
rect 31668 27004 31720 27056
rect 33048 27004 33100 27056
rect 18144 26936 18196 26988
rect 18788 26936 18840 26988
rect 20536 26979 20588 26988
rect 10968 26868 11020 26920
rect 12900 26911 12952 26920
rect 12900 26877 12909 26911
rect 12909 26877 12943 26911
rect 12943 26877 12952 26911
rect 12900 26868 12952 26877
rect 16488 26868 16540 26920
rect 20536 26945 20545 26979
rect 20545 26945 20579 26979
rect 20579 26945 20588 26979
rect 20536 26936 20588 26945
rect 21180 26936 21232 26988
rect 22100 26979 22152 26988
rect 22100 26945 22109 26979
rect 22109 26945 22143 26979
rect 22143 26945 22152 26979
rect 22100 26936 22152 26945
rect 19340 26868 19392 26920
rect 22192 26868 22244 26920
rect 22836 26868 22888 26920
rect 10232 26843 10284 26852
rect 10232 26809 10241 26843
rect 10241 26809 10275 26843
rect 10275 26809 10284 26843
rect 10232 26800 10284 26809
rect 27620 26936 27672 26988
rect 29276 26936 29328 26988
rect 33232 26979 33284 26988
rect 33232 26945 33250 26979
rect 33250 26945 33284 26979
rect 33232 26936 33284 26945
rect 34060 26936 34112 26988
rect 26240 26868 26292 26920
rect 26976 26843 27028 26852
rect 26976 26809 26985 26843
rect 26985 26809 27019 26843
rect 27019 26809 27028 26843
rect 26976 26800 27028 26809
rect 8760 26775 8812 26784
rect 8760 26741 8769 26775
rect 8769 26741 8803 26775
rect 8803 26741 8812 26775
rect 8760 26732 8812 26741
rect 14740 26775 14792 26784
rect 14740 26741 14749 26775
rect 14749 26741 14783 26775
rect 14783 26741 14792 26775
rect 14740 26732 14792 26741
rect 15200 26732 15252 26784
rect 16396 26732 16448 26784
rect 16948 26775 17000 26784
rect 16948 26741 16957 26775
rect 16957 26741 16991 26775
rect 16991 26741 17000 26775
rect 16948 26732 17000 26741
rect 17960 26732 18012 26784
rect 18328 26775 18380 26784
rect 18328 26741 18337 26775
rect 18337 26741 18371 26775
rect 18371 26741 18380 26775
rect 18328 26732 18380 26741
rect 22192 26732 22244 26784
rect 22468 26732 22520 26784
rect 22836 26775 22888 26784
rect 22836 26741 22845 26775
rect 22845 26741 22879 26775
rect 22879 26741 22888 26775
rect 22836 26732 22888 26741
rect 23204 26732 23256 26784
rect 30656 26732 30708 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 9128 26571 9180 26580
rect 9128 26537 9137 26571
rect 9137 26537 9171 26571
rect 9171 26537 9180 26571
rect 9128 26528 9180 26537
rect 11244 26571 11296 26580
rect 11244 26537 11253 26571
rect 11253 26537 11287 26571
rect 11287 26537 11296 26571
rect 11244 26528 11296 26537
rect 17132 26571 17184 26580
rect 17132 26537 17141 26571
rect 17141 26537 17175 26571
rect 17175 26537 17184 26571
rect 17132 26528 17184 26537
rect 19064 26528 19116 26580
rect 11888 26503 11940 26512
rect 9588 26392 9640 26444
rect 7380 26324 7432 26376
rect 10968 26392 11020 26444
rect 11888 26469 11897 26503
rect 11897 26469 11931 26503
rect 11931 26469 11940 26503
rect 11888 26460 11940 26469
rect 11520 26324 11572 26376
rect 11704 26367 11756 26376
rect 11704 26333 11713 26367
rect 11713 26333 11747 26367
rect 11747 26333 11756 26367
rect 11704 26324 11756 26333
rect 12256 26324 12308 26376
rect 12900 26324 12952 26376
rect 14740 26367 14792 26376
rect 14740 26333 14749 26367
rect 14749 26333 14783 26367
rect 14783 26333 14792 26367
rect 14740 26324 14792 26333
rect 16488 26324 16540 26376
rect 16948 26367 17000 26376
rect 16948 26333 16957 26367
rect 16957 26333 16991 26367
rect 16991 26333 17000 26367
rect 16948 26324 17000 26333
rect 9864 26256 9916 26308
rect 13176 26299 13228 26308
rect 13176 26265 13185 26299
rect 13185 26265 13219 26299
rect 13219 26265 13228 26299
rect 13176 26256 13228 26265
rect 17132 26256 17184 26308
rect 13820 26188 13872 26240
rect 18512 26460 18564 26512
rect 19616 26528 19668 26580
rect 19984 26528 20036 26580
rect 20444 26571 20496 26580
rect 20444 26537 20453 26571
rect 20453 26537 20487 26571
rect 20487 26537 20496 26571
rect 20444 26528 20496 26537
rect 21180 26571 21232 26580
rect 21180 26537 21189 26571
rect 21189 26537 21223 26571
rect 21223 26537 21232 26571
rect 21180 26528 21232 26537
rect 22192 26528 22244 26580
rect 29000 26528 29052 26580
rect 36636 26528 36688 26580
rect 37004 26528 37056 26580
rect 23756 26460 23808 26512
rect 33232 26460 33284 26512
rect 33416 26460 33468 26512
rect 17960 26435 18012 26444
rect 17960 26401 17969 26435
rect 17969 26401 18003 26435
rect 18003 26401 18012 26435
rect 17960 26392 18012 26401
rect 19524 26392 19576 26444
rect 20168 26392 20220 26444
rect 24308 26392 24360 26444
rect 31944 26392 31996 26444
rect 32312 26392 32364 26444
rect 33048 26392 33100 26444
rect 19248 26324 19300 26376
rect 20352 26324 20404 26376
rect 21456 26324 21508 26376
rect 27804 26367 27856 26376
rect 27804 26333 27813 26367
rect 27813 26333 27847 26367
rect 27847 26333 27856 26367
rect 27804 26324 27856 26333
rect 30380 26324 30432 26376
rect 17960 26188 18012 26240
rect 18328 26256 18380 26308
rect 19064 26256 19116 26308
rect 20076 26256 20128 26308
rect 22376 26299 22428 26308
rect 22376 26265 22385 26299
rect 22385 26265 22419 26299
rect 22419 26265 22428 26299
rect 22376 26256 22428 26265
rect 23020 26299 23072 26308
rect 23020 26265 23029 26299
rect 23029 26265 23063 26299
rect 23063 26265 23072 26299
rect 23020 26256 23072 26265
rect 26240 26299 26292 26308
rect 26240 26265 26249 26299
rect 26249 26265 26283 26299
rect 26283 26265 26292 26299
rect 26240 26256 26292 26265
rect 31484 26324 31536 26376
rect 33416 26324 33468 26376
rect 35348 26367 35400 26376
rect 35348 26333 35357 26367
rect 35357 26333 35391 26367
rect 35391 26333 35400 26367
rect 35348 26324 35400 26333
rect 33140 26256 33192 26308
rect 19616 26231 19668 26240
rect 19616 26197 19625 26231
rect 19625 26197 19659 26231
rect 19659 26197 19668 26231
rect 19616 26188 19668 26197
rect 19984 26231 20036 26240
rect 19984 26197 19993 26231
rect 19993 26197 20027 26231
rect 20027 26197 20036 26231
rect 19984 26188 20036 26197
rect 35532 26231 35584 26240
rect 35532 26197 35541 26231
rect 35541 26197 35575 26231
rect 35575 26197 35584 26231
rect 35532 26188 35584 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 9496 25984 9548 26036
rect 15844 25984 15896 26036
rect 16948 25984 17000 26036
rect 18420 25984 18472 26036
rect 19064 25984 19116 26036
rect 20536 25984 20588 26036
rect 29276 25984 29328 26036
rect 17040 25959 17092 25968
rect 17040 25925 17049 25959
rect 17049 25925 17083 25959
rect 17083 25925 17092 25959
rect 17040 25916 17092 25925
rect 23020 25916 23072 25968
rect 35532 25984 35584 26036
rect 36728 26027 36780 26036
rect 30380 25959 30432 25968
rect 30380 25925 30389 25959
rect 30389 25925 30423 25959
rect 30423 25925 30432 25959
rect 30380 25916 30432 25925
rect 32312 25916 32364 25968
rect 36728 25993 36737 26027
rect 36737 25993 36771 26027
rect 36771 25993 36780 26027
rect 36728 25984 36780 25993
rect 37832 26027 37884 26036
rect 37832 25993 37841 26027
rect 37841 25993 37875 26027
rect 37875 25993 37884 26027
rect 37832 25984 37884 25993
rect 8760 25848 8812 25900
rect 17408 25848 17460 25900
rect 17132 25823 17184 25832
rect 17132 25789 17141 25823
rect 17141 25789 17175 25823
rect 17175 25789 17184 25823
rect 17132 25780 17184 25789
rect 16488 25712 16540 25764
rect 17960 25780 18012 25832
rect 24952 25848 25004 25900
rect 25228 25891 25280 25900
rect 25228 25857 25246 25891
rect 25246 25857 25280 25891
rect 25228 25848 25280 25857
rect 33416 25848 33468 25900
rect 38016 25891 38068 25900
rect 38016 25857 38025 25891
rect 38025 25857 38059 25891
rect 38059 25857 38068 25891
rect 38016 25848 38068 25857
rect 20076 25712 20128 25764
rect 20536 25712 20588 25764
rect 22560 25780 22612 25832
rect 26240 25780 26292 25832
rect 9864 25644 9916 25696
rect 10784 25687 10836 25696
rect 10784 25653 10793 25687
rect 10793 25653 10827 25687
rect 10827 25653 10836 25687
rect 10784 25644 10836 25653
rect 12164 25644 12216 25696
rect 12348 25644 12400 25696
rect 15568 25687 15620 25696
rect 15568 25653 15577 25687
rect 15577 25653 15611 25687
rect 15611 25653 15620 25687
rect 15568 25644 15620 25653
rect 19064 25644 19116 25696
rect 20168 25644 20220 25696
rect 34612 25644 34664 25696
rect 34796 25644 34848 25696
rect 36360 25644 36412 25696
rect 36636 25644 36688 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 8576 25440 8628 25492
rect 11060 25440 11112 25492
rect 10232 25415 10284 25424
rect 8944 25304 8996 25356
rect 10232 25381 10241 25415
rect 10241 25381 10275 25415
rect 10275 25381 10284 25415
rect 10232 25372 10284 25381
rect 12164 25372 12216 25424
rect 13728 25440 13780 25492
rect 15476 25440 15528 25492
rect 18972 25440 19024 25492
rect 13452 25415 13504 25424
rect 13452 25381 13461 25415
rect 13461 25381 13495 25415
rect 13495 25381 13504 25415
rect 13452 25372 13504 25381
rect 9588 25347 9640 25356
rect 9588 25313 9597 25347
rect 9597 25313 9631 25347
rect 9631 25313 9640 25347
rect 9588 25304 9640 25313
rect 12256 25347 12308 25356
rect 12256 25313 12265 25347
rect 12265 25313 12299 25347
rect 12299 25313 12308 25347
rect 12256 25304 12308 25313
rect 12440 25304 12492 25356
rect 13452 25236 13504 25288
rect 15016 25304 15068 25356
rect 16488 25304 16540 25356
rect 17960 25304 18012 25356
rect 20168 25372 20220 25424
rect 20352 25372 20404 25424
rect 34060 25440 34112 25492
rect 35348 25483 35400 25492
rect 35348 25449 35357 25483
rect 35357 25449 35391 25483
rect 35391 25449 35400 25483
rect 35348 25440 35400 25449
rect 22652 25415 22704 25424
rect 22652 25381 22661 25415
rect 22661 25381 22695 25415
rect 22695 25381 22704 25415
rect 22652 25372 22704 25381
rect 18144 25304 18196 25356
rect 35716 25372 35768 25424
rect 29276 25304 29328 25356
rect 36360 25304 36412 25356
rect 16672 25236 16724 25288
rect 17408 25279 17460 25288
rect 17408 25245 17417 25279
rect 17417 25245 17451 25279
rect 17451 25245 17460 25279
rect 17408 25236 17460 25245
rect 18420 25236 18472 25288
rect 15568 25168 15620 25220
rect 16304 25168 16356 25220
rect 20076 25168 20128 25220
rect 20628 25236 20680 25288
rect 22468 25279 22520 25288
rect 22468 25245 22477 25279
rect 22477 25245 22511 25279
rect 22511 25245 22520 25279
rect 22468 25236 22520 25245
rect 23756 25236 23808 25288
rect 26240 25236 26292 25288
rect 29000 25236 29052 25288
rect 33692 25279 33744 25288
rect 33692 25245 33701 25279
rect 33701 25245 33735 25279
rect 33735 25245 33744 25279
rect 33692 25236 33744 25245
rect 34704 25279 34756 25288
rect 34704 25245 34713 25279
rect 34713 25245 34747 25279
rect 34747 25245 34756 25279
rect 34704 25236 34756 25245
rect 35532 25279 35584 25288
rect 35532 25245 35541 25279
rect 35541 25245 35575 25279
rect 35575 25245 35584 25279
rect 35532 25236 35584 25245
rect 35716 25279 35768 25288
rect 35716 25245 35725 25279
rect 35725 25245 35759 25279
rect 35759 25245 35768 25279
rect 35716 25236 35768 25245
rect 22192 25168 22244 25220
rect 22836 25168 22888 25220
rect 24400 25168 24452 25220
rect 26332 25168 26384 25220
rect 32312 25168 32364 25220
rect 10416 25100 10468 25152
rect 12348 25100 12400 25152
rect 14096 25143 14148 25152
rect 14096 25109 14105 25143
rect 14105 25109 14139 25143
rect 14139 25109 14148 25143
rect 14096 25100 14148 25109
rect 18052 25100 18104 25152
rect 20352 25100 20404 25152
rect 20628 25143 20680 25152
rect 20628 25109 20637 25143
rect 20637 25109 20671 25143
rect 20671 25109 20680 25143
rect 20628 25100 20680 25109
rect 20996 25100 21048 25152
rect 21824 25143 21876 25152
rect 21824 25109 21833 25143
rect 21833 25109 21867 25143
rect 21867 25109 21876 25143
rect 21824 25100 21876 25109
rect 23664 25100 23716 25152
rect 30656 25100 30708 25152
rect 30932 25143 30984 25152
rect 30932 25109 30941 25143
rect 30941 25109 30975 25143
rect 30975 25109 30984 25143
rect 30932 25100 30984 25109
rect 31024 25100 31076 25152
rect 31944 25100 31996 25152
rect 35992 25168 36044 25220
rect 37832 25100 37884 25152
rect 38200 25100 38252 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9588 24896 9640 24948
rect 10784 24896 10836 24948
rect 13636 24939 13688 24948
rect 13636 24905 13645 24939
rect 13645 24905 13679 24939
rect 13679 24905 13688 24939
rect 13636 24896 13688 24905
rect 14832 24939 14884 24948
rect 14832 24905 14841 24939
rect 14841 24905 14875 24939
rect 14875 24905 14884 24939
rect 14832 24896 14884 24905
rect 17500 24896 17552 24948
rect 20996 24896 21048 24948
rect 31024 24896 31076 24948
rect 37648 24896 37700 24948
rect 11428 24828 11480 24880
rect 17684 24828 17736 24880
rect 11980 24735 12032 24744
rect 11980 24701 11989 24735
rect 11989 24701 12023 24735
rect 12023 24701 12032 24735
rect 11980 24692 12032 24701
rect 12164 24735 12216 24744
rect 12164 24701 12173 24735
rect 12173 24701 12207 24735
rect 12207 24701 12216 24735
rect 12164 24692 12216 24701
rect 11520 24667 11572 24676
rect 11520 24633 11529 24667
rect 11529 24633 11563 24667
rect 11563 24633 11572 24667
rect 11520 24624 11572 24633
rect 13452 24692 13504 24744
rect 14096 24760 14148 24812
rect 15292 24760 15344 24812
rect 16672 24803 16724 24812
rect 16672 24769 16681 24803
rect 16681 24769 16715 24803
rect 16715 24769 16724 24803
rect 16672 24760 16724 24769
rect 19064 24803 19116 24812
rect 19064 24769 19073 24803
rect 19073 24769 19107 24803
rect 19107 24769 19116 24803
rect 19064 24760 19116 24769
rect 22192 24803 22244 24812
rect 22192 24769 22201 24803
rect 22201 24769 22235 24803
rect 22235 24769 22244 24803
rect 22192 24760 22244 24769
rect 22376 24803 22428 24812
rect 22376 24769 22385 24803
rect 22385 24769 22419 24803
rect 22419 24769 22428 24803
rect 22376 24760 22428 24769
rect 13820 24735 13872 24744
rect 13820 24701 13829 24735
rect 13829 24701 13863 24735
rect 13863 24701 13872 24735
rect 15016 24735 15068 24744
rect 13820 24692 13872 24701
rect 15016 24701 15025 24735
rect 15025 24701 15059 24735
rect 15059 24701 15068 24735
rect 15016 24692 15068 24701
rect 13268 24667 13320 24676
rect 13268 24633 13277 24667
rect 13277 24633 13311 24667
rect 13311 24633 13320 24667
rect 13268 24624 13320 24633
rect 14280 24624 14332 24676
rect 17224 24667 17276 24676
rect 17224 24633 17233 24667
rect 17233 24633 17267 24667
rect 17267 24633 17276 24667
rect 17224 24624 17276 24633
rect 17500 24692 17552 24744
rect 17960 24692 18012 24744
rect 19616 24692 19668 24744
rect 20076 24692 20128 24744
rect 20168 24735 20220 24744
rect 20168 24701 20177 24735
rect 20177 24701 20211 24735
rect 20211 24701 20220 24735
rect 20168 24692 20220 24701
rect 20628 24692 20680 24744
rect 21272 24692 21324 24744
rect 23480 24692 23532 24744
rect 20720 24624 20772 24676
rect 21180 24624 21232 24676
rect 29276 24760 29328 24812
rect 29552 24803 29604 24812
rect 29552 24769 29561 24803
rect 29561 24769 29595 24803
rect 29595 24769 29604 24803
rect 29552 24760 29604 24769
rect 31208 24803 31260 24812
rect 31208 24769 31217 24803
rect 31217 24769 31251 24803
rect 31251 24769 31260 24803
rect 31208 24760 31260 24769
rect 32128 24760 32180 24812
rect 33140 24760 33192 24812
rect 35348 24760 35400 24812
rect 29184 24692 29236 24744
rect 34520 24692 34572 24744
rect 27712 24667 27764 24676
rect 27712 24633 27721 24667
rect 27721 24633 27755 24667
rect 27755 24633 27764 24667
rect 27712 24624 27764 24633
rect 29736 24667 29788 24676
rect 29736 24633 29745 24667
rect 29745 24633 29779 24667
rect 29779 24633 29788 24667
rect 29736 24624 29788 24633
rect 31392 24667 31444 24676
rect 31392 24633 31401 24667
rect 31401 24633 31435 24667
rect 31435 24633 31444 24667
rect 31392 24624 31444 24633
rect 33232 24667 33284 24676
rect 33232 24633 33241 24667
rect 33241 24633 33275 24667
rect 33275 24633 33284 24667
rect 33232 24624 33284 24633
rect 33784 24624 33836 24676
rect 36820 24692 36872 24744
rect 35992 24624 36044 24676
rect 36176 24667 36228 24676
rect 36176 24633 36185 24667
rect 36185 24633 36219 24667
rect 36219 24633 36228 24667
rect 36176 24624 36228 24633
rect 23204 24556 23256 24608
rect 23388 24556 23440 24608
rect 23572 24556 23624 24608
rect 29828 24556 29880 24608
rect 31576 24556 31628 24608
rect 33600 24556 33652 24608
rect 34336 24599 34388 24608
rect 34336 24565 34345 24599
rect 34345 24565 34379 24599
rect 34379 24565 34388 24599
rect 37832 24624 37884 24676
rect 34336 24556 34388 24565
rect 36820 24556 36872 24608
rect 37924 24556 37976 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 13636 24352 13688 24404
rect 17684 24352 17736 24404
rect 21180 24395 21232 24404
rect 21180 24361 21189 24395
rect 21189 24361 21223 24395
rect 21223 24361 21232 24395
rect 21180 24352 21232 24361
rect 22100 24395 22152 24404
rect 22100 24361 22109 24395
rect 22109 24361 22143 24395
rect 22143 24361 22152 24395
rect 22100 24352 22152 24361
rect 23388 24352 23440 24404
rect 26424 24352 26476 24404
rect 29184 24352 29236 24404
rect 29552 24395 29604 24404
rect 29552 24361 29561 24395
rect 29561 24361 29595 24395
rect 29595 24361 29604 24395
rect 29552 24352 29604 24361
rect 32128 24395 32180 24404
rect 32128 24361 32137 24395
rect 32137 24361 32171 24395
rect 32171 24361 32180 24395
rect 32128 24352 32180 24361
rect 35440 24352 35492 24404
rect 36544 24395 36596 24404
rect 36544 24361 36553 24395
rect 36553 24361 36587 24395
rect 36587 24361 36596 24395
rect 36544 24352 36596 24361
rect 38016 24352 38068 24404
rect 16120 24284 16172 24336
rect 20076 24284 20128 24336
rect 19616 24259 19668 24268
rect 19616 24225 19625 24259
rect 19625 24225 19659 24259
rect 19659 24225 19668 24259
rect 24860 24284 24912 24336
rect 25044 24327 25096 24336
rect 25044 24293 25053 24327
rect 25053 24293 25087 24327
rect 25087 24293 25096 24327
rect 25044 24284 25096 24293
rect 19616 24216 19668 24225
rect 22836 24216 22888 24268
rect 23388 24216 23440 24268
rect 18512 24191 18564 24200
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 19892 24148 19944 24200
rect 26332 24216 26384 24268
rect 32220 24284 32272 24336
rect 33232 24216 33284 24268
rect 34152 24216 34204 24268
rect 18880 24080 18932 24132
rect 23756 24148 23808 24200
rect 28080 24148 28132 24200
rect 28908 24148 28960 24200
rect 29828 24191 29880 24200
rect 29828 24157 29837 24191
rect 29837 24157 29871 24191
rect 29871 24157 29880 24191
rect 29828 24148 29880 24157
rect 30012 24148 30064 24200
rect 31024 24191 31076 24200
rect 31024 24157 31033 24191
rect 31033 24157 31067 24191
rect 31067 24157 31076 24191
rect 31024 24148 31076 24157
rect 31576 24148 31628 24200
rect 32036 24148 32088 24200
rect 34336 24148 34388 24200
rect 34520 24148 34572 24200
rect 35716 24284 35768 24336
rect 34796 24148 34848 24200
rect 35716 24191 35768 24200
rect 35716 24157 35725 24191
rect 35725 24157 35759 24191
rect 35759 24157 35768 24191
rect 35716 24148 35768 24157
rect 21824 24080 21876 24132
rect 9128 24012 9180 24064
rect 11980 24012 12032 24064
rect 15292 24055 15344 24064
rect 15292 24021 15301 24055
rect 15301 24021 15335 24055
rect 15335 24021 15344 24055
rect 15292 24012 15344 24021
rect 17500 24012 17552 24064
rect 18696 24055 18748 24064
rect 18696 24021 18705 24055
rect 18705 24021 18739 24055
rect 18739 24021 18748 24055
rect 18696 24012 18748 24021
rect 23664 24080 23716 24132
rect 24860 24080 24912 24132
rect 30840 24080 30892 24132
rect 23388 24055 23440 24064
rect 23388 24021 23397 24055
rect 23397 24021 23431 24055
rect 23431 24021 23440 24055
rect 23388 24012 23440 24021
rect 25504 24012 25556 24064
rect 26148 24012 26200 24064
rect 34612 24080 34664 24132
rect 36452 24148 36504 24200
rect 37924 24191 37976 24200
rect 37924 24157 37933 24191
rect 37933 24157 37967 24191
rect 37967 24157 37976 24191
rect 37924 24148 37976 24157
rect 32680 24012 32732 24064
rect 33600 24012 33652 24064
rect 34152 24012 34204 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 17592 23808 17644 23860
rect 18880 23851 18932 23860
rect 18880 23817 18889 23851
rect 18889 23817 18923 23851
rect 18923 23817 18932 23851
rect 18880 23808 18932 23817
rect 19340 23808 19392 23860
rect 20076 23808 20128 23860
rect 22376 23808 22428 23860
rect 23572 23808 23624 23860
rect 23756 23851 23808 23860
rect 23756 23817 23765 23851
rect 23765 23817 23799 23851
rect 23799 23817 23808 23851
rect 23756 23808 23808 23817
rect 28356 23808 28408 23860
rect 31024 23808 31076 23860
rect 31208 23851 31260 23860
rect 31208 23817 31217 23851
rect 31217 23817 31251 23851
rect 31251 23817 31260 23851
rect 31208 23808 31260 23817
rect 33140 23808 33192 23860
rect 34796 23851 34848 23860
rect 34796 23817 34805 23851
rect 34805 23817 34839 23851
rect 34839 23817 34848 23851
rect 34796 23808 34848 23817
rect 11796 23468 11848 23520
rect 25044 23740 25096 23792
rect 25964 23783 26016 23792
rect 25964 23749 25973 23783
rect 25973 23749 26007 23783
rect 26007 23749 26016 23783
rect 25964 23740 26016 23749
rect 26608 23740 26660 23792
rect 30196 23740 30248 23792
rect 37740 23740 37792 23792
rect 18696 23715 18748 23724
rect 16948 23647 17000 23656
rect 16948 23613 16957 23647
rect 16957 23613 16991 23647
rect 16991 23613 17000 23647
rect 16948 23604 17000 23613
rect 18696 23681 18705 23715
rect 18705 23681 18739 23715
rect 18739 23681 18748 23715
rect 18696 23672 18748 23681
rect 21456 23672 21508 23724
rect 23480 23715 23532 23724
rect 23480 23681 23489 23715
rect 23489 23681 23523 23715
rect 23523 23681 23532 23715
rect 23480 23672 23532 23681
rect 24584 23715 24636 23724
rect 18788 23604 18840 23656
rect 20168 23604 20220 23656
rect 20628 23604 20680 23656
rect 22836 23647 22888 23656
rect 22836 23613 22845 23647
rect 22845 23613 22879 23647
rect 22879 23613 22888 23647
rect 22836 23604 22888 23613
rect 24584 23681 24593 23715
rect 24593 23681 24627 23715
rect 24627 23681 24636 23715
rect 24584 23672 24636 23681
rect 29552 23672 29604 23724
rect 30656 23672 30708 23724
rect 30840 23715 30892 23724
rect 30840 23681 30849 23715
rect 30849 23681 30883 23715
rect 30883 23681 30892 23715
rect 30840 23672 30892 23681
rect 31024 23715 31076 23724
rect 31024 23681 31033 23715
rect 31033 23681 31067 23715
rect 31067 23681 31076 23715
rect 31024 23672 31076 23681
rect 32680 23715 32732 23724
rect 32680 23681 32689 23715
rect 32689 23681 32723 23715
rect 32723 23681 32732 23715
rect 32680 23672 32732 23681
rect 26056 23647 26108 23656
rect 26056 23613 26065 23647
rect 26065 23613 26099 23647
rect 26099 23613 26108 23647
rect 26056 23604 26108 23613
rect 26148 23647 26200 23656
rect 26148 23613 26157 23647
rect 26157 23613 26191 23647
rect 26191 23613 26200 23647
rect 26148 23604 26200 23613
rect 29644 23647 29696 23656
rect 29644 23613 29653 23647
rect 29653 23613 29687 23647
rect 29687 23613 29696 23647
rect 29644 23604 29696 23613
rect 32496 23647 32548 23656
rect 32496 23613 32505 23647
rect 32505 23613 32539 23647
rect 32539 23613 32548 23647
rect 34520 23672 34572 23724
rect 32496 23604 32548 23613
rect 34152 23647 34204 23656
rect 34152 23613 34161 23647
rect 34161 23613 34195 23647
rect 34195 23613 34204 23647
rect 34152 23604 34204 23613
rect 19064 23468 19116 23520
rect 23020 23536 23072 23588
rect 24676 23536 24728 23588
rect 21180 23511 21232 23520
rect 21180 23477 21189 23511
rect 21189 23477 21223 23511
rect 21223 23477 21232 23511
rect 21180 23468 21232 23477
rect 28264 23468 28316 23520
rect 37096 23468 37148 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 16948 23264 17000 23316
rect 17408 23264 17460 23316
rect 22008 23264 22060 23316
rect 24584 23264 24636 23316
rect 26608 23307 26660 23316
rect 26608 23273 26617 23307
rect 26617 23273 26651 23307
rect 26651 23273 26660 23307
rect 26608 23264 26660 23273
rect 29276 23264 29328 23316
rect 29552 23307 29604 23316
rect 29552 23273 29561 23307
rect 29561 23273 29595 23307
rect 29595 23273 29604 23307
rect 29552 23264 29604 23273
rect 30196 23307 30248 23316
rect 30196 23273 30205 23307
rect 30205 23273 30239 23307
rect 30239 23273 30248 23307
rect 30196 23264 30248 23273
rect 31760 23307 31812 23316
rect 31760 23273 31769 23307
rect 31769 23273 31803 23307
rect 31803 23273 31812 23307
rect 31760 23264 31812 23273
rect 32496 23307 32548 23316
rect 32496 23273 32505 23307
rect 32505 23273 32539 23307
rect 32539 23273 32548 23307
rect 32496 23264 32548 23273
rect 34704 23307 34756 23316
rect 34704 23273 34713 23307
rect 34713 23273 34747 23307
rect 34747 23273 34756 23307
rect 34704 23264 34756 23273
rect 35716 23264 35768 23316
rect 35900 23264 35952 23316
rect 20352 23196 20404 23248
rect 20628 23128 20680 23180
rect 25872 23128 25924 23180
rect 23020 23103 23072 23112
rect 23020 23069 23029 23103
rect 23029 23069 23063 23103
rect 23063 23069 23072 23103
rect 23020 23060 23072 23069
rect 23848 23060 23900 23112
rect 20812 22992 20864 23044
rect 21180 22992 21232 23044
rect 21732 22967 21784 22976
rect 21732 22933 21741 22967
rect 21741 22933 21775 22967
rect 21775 22933 21784 22967
rect 22836 22992 22888 23044
rect 24676 23060 24728 23112
rect 25228 23103 25280 23112
rect 25228 23069 25237 23103
rect 25237 23069 25271 23103
rect 25271 23069 25280 23103
rect 25228 23060 25280 23069
rect 29644 23128 29696 23180
rect 35348 23196 35400 23248
rect 34152 23128 34204 23180
rect 34520 23128 34572 23180
rect 28264 23103 28316 23112
rect 28264 23069 28273 23103
rect 28273 23069 28307 23103
rect 28307 23069 28316 23103
rect 28264 23060 28316 23069
rect 30380 23060 30432 23112
rect 30932 23103 30984 23112
rect 30932 23069 30941 23103
rect 30941 23069 30975 23103
rect 30975 23069 30984 23103
rect 30932 23060 30984 23069
rect 32496 23060 32548 23112
rect 33140 23103 33192 23112
rect 33140 23069 33149 23103
rect 33149 23069 33183 23103
rect 33183 23069 33192 23103
rect 33140 23060 33192 23069
rect 34888 23103 34940 23112
rect 34888 23069 34897 23103
rect 34897 23069 34931 23103
rect 34931 23069 34940 23103
rect 34888 23060 34940 23069
rect 37004 23103 37056 23112
rect 23112 22967 23164 22976
rect 21732 22924 21784 22933
rect 23112 22933 23121 22967
rect 23121 22933 23155 22967
rect 23155 22933 23164 22967
rect 23112 22924 23164 22933
rect 24400 22924 24452 22976
rect 31852 22992 31904 23044
rect 37004 23069 37013 23103
rect 37013 23069 37047 23103
rect 37047 23069 37056 23103
rect 37004 23060 37056 23069
rect 27712 22924 27764 22976
rect 35900 22924 35952 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 23112 22720 23164 22772
rect 25228 22720 25280 22772
rect 30012 22763 30064 22772
rect 23848 22695 23900 22704
rect 20628 22584 20680 22636
rect 21824 22584 21876 22636
rect 22560 22584 22612 22636
rect 21732 22516 21784 22568
rect 22100 22559 22152 22568
rect 22100 22525 22109 22559
rect 22109 22525 22143 22559
rect 22143 22525 22152 22559
rect 22100 22516 22152 22525
rect 23848 22661 23857 22695
rect 23857 22661 23891 22695
rect 23891 22661 23900 22695
rect 23848 22652 23900 22661
rect 24400 22695 24452 22704
rect 24400 22661 24409 22695
rect 24409 22661 24443 22695
rect 24443 22661 24452 22695
rect 24400 22652 24452 22661
rect 30012 22729 30021 22763
rect 30021 22729 30055 22763
rect 30055 22729 30064 22763
rect 30012 22720 30064 22729
rect 30840 22720 30892 22772
rect 32312 22763 32364 22772
rect 32312 22729 32321 22763
rect 32321 22729 32355 22763
rect 32355 22729 32364 22763
rect 32312 22720 32364 22729
rect 32496 22720 32548 22772
rect 30564 22652 30616 22704
rect 25596 22627 25648 22636
rect 25596 22593 25605 22627
rect 25605 22593 25639 22627
rect 25639 22593 25648 22627
rect 25596 22584 25648 22593
rect 27712 22627 27764 22636
rect 27712 22593 27721 22627
rect 27721 22593 27755 22627
rect 27755 22593 27764 22627
rect 27712 22584 27764 22593
rect 28356 22627 28408 22636
rect 28356 22593 28365 22627
rect 28365 22593 28399 22627
rect 28399 22593 28408 22627
rect 28356 22584 28408 22593
rect 29828 22627 29880 22636
rect 29828 22593 29837 22627
rect 29837 22593 29871 22627
rect 29871 22593 29880 22627
rect 29828 22584 29880 22593
rect 30196 22584 30248 22636
rect 27620 22516 27672 22568
rect 30380 22516 30432 22568
rect 33692 22720 33744 22772
rect 34888 22720 34940 22772
rect 36360 22720 36412 22772
rect 35716 22695 35768 22704
rect 35716 22661 35725 22695
rect 35725 22661 35759 22695
rect 35759 22661 35768 22695
rect 35716 22652 35768 22661
rect 34704 22584 34756 22636
rect 35808 22559 35860 22568
rect 35808 22525 35817 22559
rect 35817 22525 35851 22559
rect 35851 22525 35860 22559
rect 35808 22516 35860 22525
rect 30472 22448 30524 22500
rect 30748 22448 30800 22500
rect 34612 22380 34664 22432
rect 38108 22380 38160 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 25596 22176 25648 22228
rect 28356 22176 28408 22228
rect 33140 22176 33192 22228
rect 34704 22219 34756 22228
rect 34704 22185 34713 22219
rect 34713 22185 34747 22219
rect 34747 22185 34756 22219
rect 34704 22176 34756 22185
rect 35900 22219 35952 22228
rect 35900 22185 35909 22219
rect 35909 22185 35943 22219
rect 35943 22185 35952 22219
rect 35900 22176 35952 22185
rect 10968 22108 11020 22160
rect 11980 22108 12032 22160
rect 22560 22108 22612 22160
rect 28172 22108 28224 22160
rect 25504 22040 25556 22092
rect 26792 22083 26844 22092
rect 26792 22049 26801 22083
rect 26801 22049 26835 22083
rect 26835 22049 26844 22083
rect 26792 22040 26844 22049
rect 27620 22083 27672 22092
rect 27620 22049 27629 22083
rect 27629 22049 27663 22083
rect 27663 22049 27672 22083
rect 30380 22108 30432 22160
rect 31484 22108 31536 22160
rect 27620 22040 27672 22049
rect 30196 22083 30248 22092
rect 30196 22049 30205 22083
rect 30205 22049 30239 22083
rect 30239 22049 30248 22083
rect 30196 22040 30248 22049
rect 30288 22040 30340 22092
rect 35808 22040 35860 22092
rect 16396 21972 16448 22024
rect 20352 21972 20404 22024
rect 21824 22015 21876 22024
rect 21824 21981 21833 22015
rect 21833 21981 21867 22015
rect 21867 21981 21876 22015
rect 21824 21972 21876 21981
rect 22100 21972 22152 22024
rect 26976 21972 27028 22024
rect 27988 21972 28040 22024
rect 28632 22015 28684 22024
rect 28632 21981 28641 22015
rect 28641 21981 28675 22015
rect 28675 21981 28684 22015
rect 28632 21972 28684 21981
rect 30012 22015 30064 22024
rect 30012 21981 30021 22015
rect 30021 21981 30055 22015
rect 30055 21981 30064 22015
rect 30012 21972 30064 21981
rect 34612 21972 34664 22024
rect 35624 21972 35676 22024
rect 36268 22015 36320 22024
rect 36268 21981 36277 22015
rect 36277 21981 36311 22015
rect 36311 21981 36320 22015
rect 36268 21972 36320 21981
rect 27252 21904 27304 21956
rect 30104 21904 30156 21956
rect 22100 21879 22152 21888
rect 22100 21845 22109 21879
rect 22109 21845 22143 21879
rect 22143 21845 22152 21879
rect 22100 21836 22152 21845
rect 27160 21836 27212 21888
rect 28080 21836 28132 21888
rect 32772 21836 32824 21888
rect 35440 21836 35492 21888
rect 37372 21836 37424 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 28632 21675 28684 21684
rect 28632 21641 28641 21675
rect 28641 21641 28675 21675
rect 28675 21641 28684 21675
rect 28632 21632 28684 21641
rect 31024 21632 31076 21684
rect 34796 21632 34848 21684
rect 37004 21632 37056 21684
rect 31392 21564 31444 21616
rect 32864 21496 32916 21548
rect 36268 21539 36320 21548
rect 36268 21505 36277 21539
rect 36277 21505 36311 21539
rect 36311 21505 36320 21539
rect 36268 21496 36320 21505
rect 26792 21428 26844 21480
rect 27160 21292 27212 21344
rect 30196 21428 30248 21480
rect 31484 21428 31536 21480
rect 36452 21428 36504 21480
rect 29368 21292 29420 21344
rect 29644 21335 29696 21344
rect 29644 21301 29653 21335
rect 29653 21301 29687 21335
rect 29687 21301 29696 21335
rect 29644 21292 29696 21301
rect 32772 21292 32824 21344
rect 35440 21292 35492 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 27252 21131 27304 21140
rect 27252 21097 27261 21131
rect 27261 21097 27295 21131
rect 27295 21097 27304 21131
rect 27252 21088 27304 21097
rect 27988 21131 28040 21140
rect 27988 21097 27997 21131
rect 27997 21097 28031 21131
rect 28031 21097 28040 21131
rect 27988 21088 28040 21097
rect 30012 21088 30064 21140
rect 30932 21131 30984 21140
rect 30932 21097 30941 21131
rect 30941 21097 30975 21131
rect 30975 21097 30984 21131
rect 30932 21088 30984 21097
rect 35532 21088 35584 21140
rect 36728 21088 36780 21140
rect 29368 21020 29420 21072
rect 35900 21020 35952 21072
rect 36820 21020 36872 21072
rect 22100 20952 22152 21004
rect 30196 20952 30248 21004
rect 35808 20952 35860 21004
rect 29460 20884 29512 20936
rect 30104 20927 30156 20936
rect 30104 20893 30113 20927
rect 30113 20893 30147 20927
rect 30147 20893 30156 20927
rect 30104 20884 30156 20893
rect 31300 20927 31352 20936
rect 31300 20893 31309 20927
rect 31309 20893 31343 20927
rect 31343 20893 31352 20927
rect 31300 20884 31352 20893
rect 36728 20884 36780 20936
rect 28356 20859 28408 20868
rect 28356 20825 28365 20859
rect 28365 20825 28399 20859
rect 28399 20825 28408 20859
rect 28356 20816 28408 20825
rect 31668 20816 31720 20868
rect 35808 20816 35860 20868
rect 20996 20791 21048 20800
rect 20996 20757 21005 20791
rect 21005 20757 21039 20791
rect 21039 20757 21048 20791
rect 20996 20748 21048 20757
rect 28816 20748 28868 20800
rect 30748 20748 30800 20800
rect 32312 20748 32364 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 20996 20544 21048 20596
rect 27068 20544 27120 20596
rect 28356 20587 28408 20596
rect 28356 20553 28365 20587
rect 28365 20553 28399 20587
rect 28399 20553 28408 20587
rect 28356 20544 28408 20553
rect 29828 20544 29880 20596
rect 30104 20544 30156 20596
rect 23296 20476 23348 20528
rect 29920 20451 29972 20460
rect 29920 20417 29929 20451
rect 29929 20417 29963 20451
rect 29963 20417 29972 20451
rect 29920 20408 29972 20417
rect 22100 20340 22152 20392
rect 30012 20383 30064 20392
rect 30012 20349 30021 20383
rect 30021 20349 30055 20383
rect 30055 20349 30064 20383
rect 30012 20340 30064 20349
rect 30196 20383 30248 20392
rect 30196 20349 30205 20383
rect 30205 20349 30239 20383
rect 30239 20349 30248 20383
rect 30196 20340 30248 20349
rect 20168 20204 20220 20256
rect 28816 20247 28868 20256
rect 28816 20213 28825 20247
rect 28825 20213 28859 20247
rect 28859 20213 28868 20247
rect 28816 20204 28868 20213
rect 30748 20247 30800 20256
rect 30748 20213 30757 20247
rect 30757 20213 30791 20247
rect 30791 20213 30800 20247
rect 30748 20204 30800 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 21180 20000 21232 20052
rect 21364 20000 21416 20052
rect 20444 19907 20496 19916
rect 20444 19873 20453 19907
rect 20453 19873 20487 19907
rect 20487 19873 20496 19907
rect 20444 19864 20496 19873
rect 22100 19864 22152 19916
rect 22928 20000 22980 20052
rect 29184 20000 29236 20052
rect 29920 20000 29972 20052
rect 32220 20000 32272 20052
rect 36268 20000 36320 20052
rect 35900 19864 35952 19916
rect 29920 19796 29972 19848
rect 36452 19839 36504 19848
rect 36452 19805 36461 19839
rect 36461 19805 36495 19839
rect 36495 19805 36504 19839
rect 36452 19796 36504 19805
rect 30564 19728 30616 19780
rect 20076 19660 20128 19712
rect 21180 19660 21232 19712
rect 21364 19703 21416 19712
rect 21364 19669 21373 19703
rect 21373 19669 21407 19703
rect 21407 19669 21416 19703
rect 21364 19660 21416 19669
rect 22008 19660 22060 19712
rect 30104 19660 30156 19712
rect 37464 19660 37516 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 20444 19499 20496 19508
rect 20444 19465 20453 19499
rect 20453 19465 20487 19499
rect 20487 19465 20496 19499
rect 20444 19456 20496 19465
rect 21364 19456 21416 19508
rect 21824 19499 21876 19508
rect 21824 19465 21833 19499
rect 21833 19465 21867 19499
rect 21867 19465 21876 19499
rect 21824 19456 21876 19465
rect 32680 19456 32732 19508
rect 30656 19388 30708 19440
rect 36084 19456 36136 19508
rect 22100 19320 22152 19372
rect 30104 19363 30156 19372
rect 30104 19329 30113 19363
rect 30113 19329 30147 19363
rect 30147 19329 30156 19363
rect 30104 19320 30156 19329
rect 21180 19295 21232 19304
rect 21180 19261 21189 19295
rect 21189 19261 21223 19295
rect 21223 19261 21232 19295
rect 21180 19252 21232 19261
rect 27160 19252 27212 19304
rect 33508 19252 33560 19304
rect 21824 19116 21876 19168
rect 29184 19116 29236 19168
rect 29920 19116 29972 19168
rect 35900 19320 35952 19372
rect 36544 19252 36596 19304
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 22100 18776 22152 18828
rect 23388 18776 23440 18828
rect 25412 18912 25464 18964
rect 36084 18912 36136 18964
rect 26240 18640 26292 18692
rect 20720 18572 20772 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 21088 18368 21140 18420
rect 33784 18411 33836 18420
rect 33784 18377 33793 18411
rect 33793 18377 33827 18411
rect 33827 18377 33836 18411
rect 33784 18368 33836 18377
rect 16488 18232 16540 18284
rect 20444 18164 20496 18216
rect 34612 18164 34664 18216
rect 15936 18028 15988 18080
rect 33232 18028 33284 18080
rect 34796 18028 34848 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 34612 17824 34664 17876
rect 16488 17484 16540 17536
rect 34612 17484 34664 17536
rect 37740 17484 37792 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 16948 17280 17000 17332
rect 17500 17280 17552 17332
rect 18420 17280 18472 17332
rect 21548 17280 21600 17332
rect 25136 17076 25188 17128
rect 18328 17008 18380 17060
rect 33968 17280 34020 17332
rect 26424 17008 26476 17060
rect 29736 17008 29788 17060
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 24400 16736 24452 16788
rect 18420 16643 18472 16652
rect 18420 16609 18429 16643
rect 18429 16609 18463 16643
rect 18463 16609 18472 16643
rect 18420 16600 18472 16609
rect 18972 16600 19024 16652
rect 20444 16600 20496 16652
rect 23388 16532 23440 16584
rect 25136 16532 25188 16584
rect 19340 16464 19392 16516
rect 22744 16464 22796 16516
rect 16856 16396 16908 16448
rect 18328 16439 18380 16448
rect 18328 16405 18337 16439
rect 18337 16405 18371 16439
rect 18371 16405 18380 16439
rect 18328 16396 18380 16405
rect 18512 16396 18564 16448
rect 21824 16396 21876 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 17960 16192 18012 16244
rect 18604 16192 18656 16244
rect 19340 16192 19392 16244
rect 19432 16124 19484 16176
rect 24032 16124 24084 16176
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 24860 16056 24912 16108
rect 18972 16031 19024 16040
rect 18972 15997 18981 16031
rect 18981 15997 19015 16031
rect 19015 15997 19024 16031
rect 18972 15988 19024 15997
rect 22652 15988 22704 16040
rect 23296 16031 23348 16040
rect 23296 15997 23305 16031
rect 23305 15997 23339 16031
rect 23339 15997 23348 16031
rect 23296 15988 23348 15997
rect 19432 15852 19484 15904
rect 21732 15852 21784 15904
rect 22560 15852 22612 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 17960 15580 18012 15632
rect 18972 15512 19024 15564
rect 22192 15648 22244 15700
rect 30656 15648 30708 15700
rect 25596 15580 25648 15632
rect 26424 15580 26476 15632
rect 23296 15512 23348 15564
rect 17408 15444 17460 15496
rect 20352 15444 20404 15496
rect 21732 15487 21784 15496
rect 21732 15453 21741 15487
rect 21741 15453 21775 15487
rect 21775 15453 21784 15487
rect 21732 15444 21784 15453
rect 22560 15487 22612 15496
rect 17500 15376 17552 15428
rect 22560 15453 22569 15487
rect 22569 15453 22603 15487
rect 22603 15453 22612 15487
rect 22560 15444 22612 15453
rect 24400 15487 24452 15496
rect 24400 15453 24409 15487
rect 24409 15453 24443 15487
rect 24443 15453 24452 15487
rect 24400 15444 24452 15453
rect 26056 15444 26108 15496
rect 30288 15580 30340 15632
rect 36268 15512 36320 15564
rect 26608 15444 26660 15496
rect 22652 15376 22704 15428
rect 32128 15444 32180 15496
rect 33140 15444 33192 15496
rect 15476 15308 15528 15360
rect 19248 15308 19300 15360
rect 19984 15351 20036 15360
rect 19984 15317 19993 15351
rect 19993 15317 20027 15351
rect 20027 15317 20036 15351
rect 19984 15308 20036 15317
rect 20904 15308 20956 15360
rect 25412 15351 25464 15360
rect 25412 15317 25421 15351
rect 25421 15317 25455 15351
rect 25455 15317 25464 15351
rect 25412 15308 25464 15317
rect 25504 15308 25556 15360
rect 26516 15308 26568 15360
rect 33324 15376 33376 15428
rect 27528 15308 27580 15360
rect 36452 15308 36504 15360
rect 36912 15351 36964 15360
rect 36912 15317 36921 15351
rect 36921 15317 36955 15351
rect 36955 15317 36964 15351
rect 36912 15308 36964 15317
rect 37372 15308 37424 15360
rect 37924 15351 37976 15360
rect 37924 15317 37933 15351
rect 37933 15317 37967 15351
rect 37967 15317 37976 15351
rect 37924 15308 37976 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 17316 15104 17368 15156
rect 20260 15104 20312 15156
rect 20352 15104 20404 15156
rect 24400 15104 24452 15156
rect 24952 15147 25004 15156
rect 24952 15113 24961 15147
rect 24961 15113 24995 15147
rect 24995 15113 25004 15147
rect 24952 15104 25004 15113
rect 33140 15104 33192 15156
rect 20628 15036 20680 15088
rect 21640 15036 21692 15088
rect 25412 15036 25464 15088
rect 20996 14968 21048 15020
rect 22192 15011 22244 15020
rect 22192 14977 22201 15011
rect 22201 14977 22235 15011
rect 22235 14977 22244 15011
rect 22192 14968 22244 14977
rect 18972 14900 19024 14952
rect 22652 14900 22704 14952
rect 20904 14875 20956 14884
rect 20904 14841 20913 14875
rect 20913 14841 20947 14875
rect 20947 14841 20956 14875
rect 20904 14832 20956 14841
rect 17224 14807 17276 14816
rect 17224 14773 17233 14807
rect 17233 14773 17267 14807
rect 17267 14773 17276 14807
rect 17224 14764 17276 14773
rect 17408 14764 17460 14816
rect 18972 14764 19024 14816
rect 23572 14764 23624 14816
rect 25320 14968 25372 15020
rect 30288 15011 30340 15020
rect 30288 14977 30297 15011
rect 30297 14977 30331 15011
rect 30331 14977 30340 15011
rect 30288 14968 30340 14977
rect 32128 15011 32180 15020
rect 32128 14977 32137 15011
rect 32137 14977 32171 15011
rect 32171 14977 32180 15011
rect 32128 14968 32180 14977
rect 25136 14943 25188 14952
rect 25136 14909 25145 14943
rect 25145 14909 25179 14943
rect 25179 14909 25188 14943
rect 25136 14900 25188 14909
rect 25504 14900 25556 14952
rect 26056 14943 26108 14952
rect 26056 14909 26065 14943
rect 26065 14909 26099 14943
rect 26099 14909 26108 14943
rect 26056 14900 26108 14909
rect 29920 14832 29972 14884
rect 30196 14832 30248 14884
rect 28540 14764 28592 14816
rect 30472 14807 30524 14816
rect 30472 14773 30481 14807
rect 30481 14773 30515 14807
rect 30515 14773 30524 14807
rect 30472 14764 30524 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19156 14560 19208 14612
rect 20628 14560 20680 14612
rect 20996 14603 21048 14612
rect 20996 14569 21005 14603
rect 21005 14569 21039 14603
rect 21039 14569 21048 14603
rect 20996 14560 21048 14569
rect 21640 14560 21692 14612
rect 25320 14603 25372 14612
rect 25320 14569 25329 14603
rect 25329 14569 25363 14603
rect 25363 14569 25372 14603
rect 25320 14560 25372 14569
rect 26424 14603 26476 14612
rect 26424 14569 26433 14603
rect 26433 14569 26467 14603
rect 26467 14569 26476 14603
rect 26424 14560 26476 14569
rect 24952 14492 25004 14544
rect 18880 14424 18932 14476
rect 25136 14424 25188 14476
rect 25412 14424 25464 14476
rect 33692 14424 33744 14476
rect 36268 14467 36320 14476
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 17040 14356 17092 14408
rect 26608 14356 26660 14408
rect 28540 14399 28592 14408
rect 28540 14365 28549 14399
rect 28549 14365 28583 14399
rect 28583 14365 28592 14399
rect 28540 14356 28592 14365
rect 15844 14288 15896 14340
rect 17224 14288 17276 14340
rect 19340 14288 19392 14340
rect 26424 14288 26476 14340
rect 32588 14399 32640 14408
rect 32588 14365 32597 14399
rect 32597 14365 32631 14399
rect 32631 14365 32640 14399
rect 32588 14356 32640 14365
rect 15660 14263 15712 14272
rect 15660 14229 15669 14263
rect 15669 14229 15703 14263
rect 15703 14229 15712 14263
rect 15660 14220 15712 14229
rect 16580 14263 16632 14272
rect 16580 14229 16589 14263
rect 16589 14229 16623 14263
rect 16623 14229 16632 14263
rect 16580 14220 16632 14229
rect 17316 14220 17368 14272
rect 17776 14263 17828 14272
rect 17776 14229 17785 14263
rect 17785 14229 17819 14263
rect 17819 14229 17828 14263
rect 17776 14220 17828 14229
rect 18144 14263 18196 14272
rect 18144 14229 18153 14263
rect 18153 14229 18187 14263
rect 18187 14229 18196 14263
rect 18144 14220 18196 14229
rect 19156 14220 19208 14272
rect 25412 14220 25464 14272
rect 30288 14220 30340 14272
rect 31852 14263 31904 14272
rect 31852 14229 31861 14263
rect 31861 14229 31895 14263
rect 31895 14229 31904 14263
rect 31852 14220 31904 14229
rect 33416 14263 33468 14272
rect 33416 14229 33425 14263
rect 33425 14229 33459 14263
rect 33459 14229 33468 14263
rect 33416 14220 33468 14229
rect 34612 14220 34664 14272
rect 36268 14433 36277 14467
rect 36277 14433 36311 14467
rect 36311 14433 36320 14467
rect 36268 14424 36320 14433
rect 36544 14424 36596 14476
rect 36544 14263 36596 14272
rect 36544 14229 36553 14263
rect 36553 14229 36587 14263
rect 36587 14229 36596 14263
rect 36544 14220 36596 14229
rect 37280 14220 37332 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 17040 14016 17092 14068
rect 18144 14016 18196 14068
rect 18696 14059 18748 14068
rect 18696 14025 18705 14059
rect 18705 14025 18739 14059
rect 18739 14025 18748 14059
rect 18696 14016 18748 14025
rect 23756 14016 23808 14068
rect 25412 14059 25464 14068
rect 25412 14025 25421 14059
rect 25421 14025 25455 14059
rect 25455 14025 25464 14059
rect 25412 14016 25464 14025
rect 25504 14016 25556 14068
rect 31852 14016 31904 14068
rect 20996 13948 21048 14000
rect 27436 13948 27488 14000
rect 15660 13880 15712 13932
rect 18512 13880 18564 13932
rect 20168 13923 20220 13932
rect 20168 13889 20177 13923
rect 20177 13889 20211 13923
rect 20211 13889 20220 13923
rect 20168 13880 20220 13889
rect 21088 13880 21140 13932
rect 22652 13880 22704 13932
rect 25412 13880 25464 13932
rect 30104 13880 30156 13932
rect 36452 13923 36504 13932
rect 36452 13889 36461 13923
rect 36461 13889 36495 13923
rect 36495 13889 36504 13923
rect 36452 13880 36504 13889
rect 15844 13855 15896 13864
rect 15844 13821 15853 13855
rect 15853 13821 15887 13855
rect 15887 13821 15896 13855
rect 15844 13812 15896 13821
rect 17408 13812 17460 13864
rect 18236 13812 18288 13864
rect 20260 13812 20312 13864
rect 25504 13812 25556 13864
rect 20996 13744 21048 13796
rect 22192 13744 22244 13796
rect 23756 13744 23808 13796
rect 30380 13744 30432 13796
rect 19892 13676 19944 13728
rect 36268 13719 36320 13728
rect 36268 13685 36277 13719
rect 36277 13685 36311 13719
rect 36311 13685 36320 13719
rect 36268 13676 36320 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 18052 13404 18104 13456
rect 24492 13447 24544 13456
rect 24492 13413 24501 13447
rect 24501 13413 24535 13447
rect 24535 13413 24544 13447
rect 24492 13404 24544 13413
rect 14372 13311 14424 13320
rect 14372 13277 14381 13311
rect 14381 13277 14415 13311
rect 14415 13277 14424 13311
rect 14372 13268 14424 13277
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 17776 13268 17828 13320
rect 18236 13311 18288 13320
rect 18236 13277 18245 13311
rect 18245 13277 18279 13311
rect 18279 13277 18288 13311
rect 18236 13268 18288 13277
rect 19248 13311 19300 13320
rect 19248 13277 19257 13311
rect 19257 13277 19291 13311
rect 19291 13277 19300 13311
rect 19248 13268 19300 13277
rect 19892 13311 19944 13320
rect 19892 13277 19901 13311
rect 19901 13277 19935 13311
rect 19935 13277 19944 13311
rect 19892 13268 19944 13277
rect 23020 13311 23072 13320
rect 23020 13277 23029 13311
rect 23029 13277 23063 13311
rect 23063 13277 23072 13311
rect 23020 13268 23072 13277
rect 25872 13311 25924 13320
rect 25872 13277 25881 13311
rect 25881 13277 25915 13311
rect 25915 13277 25924 13311
rect 25872 13268 25924 13277
rect 22928 13200 22980 13252
rect 36636 13472 36688 13524
rect 27160 13268 27212 13320
rect 31760 13268 31812 13320
rect 38108 13311 38160 13320
rect 38108 13277 38117 13311
rect 38117 13277 38151 13311
rect 38151 13277 38160 13311
rect 38108 13268 38160 13277
rect 30288 13200 30340 13252
rect 37464 13200 37516 13252
rect 14556 13175 14608 13184
rect 14556 13141 14565 13175
rect 14565 13141 14599 13175
rect 14599 13141 14608 13175
rect 14556 13132 14608 13141
rect 17316 13132 17368 13184
rect 17408 13132 17460 13184
rect 17776 13132 17828 13184
rect 18236 13132 18288 13184
rect 18420 13175 18472 13184
rect 18420 13141 18429 13175
rect 18429 13141 18463 13175
rect 18463 13141 18472 13175
rect 18420 13132 18472 13141
rect 20076 13175 20128 13184
rect 20076 13141 20085 13175
rect 20085 13141 20119 13175
rect 20119 13141 20128 13175
rect 20076 13132 20128 13141
rect 22192 13132 22244 13184
rect 30104 13132 30156 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 14556 12928 14608 12980
rect 22928 12928 22980 12980
rect 32128 12971 32180 12980
rect 32128 12937 32137 12971
rect 32137 12937 32171 12971
rect 32171 12937 32180 12971
rect 32128 12928 32180 12937
rect 33784 12928 33836 12980
rect 37464 12971 37516 12980
rect 37464 12937 37473 12971
rect 37473 12937 37507 12971
rect 37507 12937 37516 12971
rect 37464 12928 37516 12937
rect 15936 12835 15988 12844
rect 15936 12801 15945 12835
rect 15945 12801 15979 12835
rect 15979 12801 15988 12835
rect 15936 12792 15988 12801
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 18420 12860 18472 12912
rect 18972 12835 19024 12844
rect 18972 12801 18981 12835
rect 18981 12801 19015 12835
rect 19015 12801 19024 12835
rect 18972 12792 19024 12801
rect 19984 12792 20036 12844
rect 20720 12792 20772 12844
rect 20904 12792 20956 12844
rect 23756 12792 23808 12844
rect 25504 12792 25556 12844
rect 25872 12792 25924 12844
rect 27160 12860 27212 12912
rect 29552 12860 29604 12912
rect 33416 12860 33468 12912
rect 34796 12792 34848 12844
rect 35348 12835 35400 12844
rect 35348 12801 35357 12835
rect 35357 12801 35391 12835
rect 35391 12801 35400 12835
rect 35348 12792 35400 12801
rect 37280 12835 37332 12844
rect 37280 12801 37289 12835
rect 37289 12801 37323 12835
rect 37323 12801 37332 12835
rect 37280 12792 37332 12801
rect 16672 12767 16724 12776
rect 16672 12733 16681 12767
rect 16681 12733 16715 12767
rect 16715 12733 16724 12767
rect 16672 12724 16724 12733
rect 17776 12724 17828 12776
rect 18788 12767 18840 12776
rect 18788 12733 18797 12767
rect 18797 12733 18831 12767
rect 18831 12733 18840 12767
rect 18788 12724 18840 12733
rect 19892 12724 19944 12776
rect 21088 12724 21140 12776
rect 21180 12724 21232 12776
rect 21824 12724 21876 12776
rect 23204 12767 23256 12776
rect 20628 12656 20680 12708
rect 23204 12733 23213 12767
rect 23213 12733 23247 12767
rect 23247 12733 23256 12767
rect 23204 12724 23256 12733
rect 31760 12724 31812 12776
rect 17224 12588 17276 12640
rect 19248 12588 19300 12640
rect 20076 12588 20128 12640
rect 20444 12631 20496 12640
rect 20444 12597 20453 12631
rect 20453 12597 20487 12631
rect 20487 12597 20496 12631
rect 20444 12588 20496 12597
rect 21824 12631 21876 12640
rect 21824 12597 21833 12631
rect 21833 12597 21867 12631
rect 21867 12597 21876 12631
rect 21824 12588 21876 12597
rect 23664 12631 23716 12640
rect 23664 12597 23673 12631
rect 23673 12597 23707 12631
rect 23707 12597 23716 12631
rect 23664 12588 23716 12597
rect 27252 12656 27304 12708
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 13176 12384 13228 12436
rect 13728 12384 13780 12436
rect 18236 12384 18288 12436
rect 18788 12384 18840 12436
rect 20260 12384 20312 12436
rect 21640 12427 21692 12436
rect 21640 12393 21649 12427
rect 21649 12393 21683 12427
rect 21683 12393 21692 12427
rect 21640 12384 21692 12393
rect 17500 12316 17552 12368
rect 17776 12316 17828 12368
rect 37372 12384 37424 12436
rect 16580 12180 16632 12232
rect 17960 12248 18012 12300
rect 17500 12223 17552 12232
rect 17500 12189 17509 12223
rect 17509 12189 17543 12223
rect 17543 12189 17552 12223
rect 17500 12180 17552 12189
rect 18144 12223 18196 12232
rect 18144 12189 18153 12223
rect 18153 12189 18187 12223
rect 18187 12189 18196 12223
rect 18144 12180 18196 12189
rect 19340 12180 19392 12232
rect 20260 12248 20312 12300
rect 27160 12291 27212 12300
rect 27160 12257 27169 12291
rect 27169 12257 27203 12291
rect 27203 12257 27212 12291
rect 27160 12248 27212 12257
rect 23020 12223 23072 12232
rect 23020 12189 23029 12223
rect 23029 12189 23063 12223
rect 23063 12189 23072 12223
rect 23020 12180 23072 12189
rect 23204 12180 23256 12232
rect 26608 12180 26660 12232
rect 30472 12180 30524 12232
rect 31760 12180 31812 12232
rect 31944 12180 31996 12232
rect 35348 12180 35400 12232
rect 38108 12180 38160 12232
rect 16672 12112 16724 12164
rect 16856 12112 16908 12164
rect 16580 12044 16632 12096
rect 25228 12112 25280 12164
rect 27712 12112 27764 12164
rect 36360 12155 36412 12164
rect 36360 12121 36394 12155
rect 36394 12121 36412 12155
rect 36360 12112 36412 12121
rect 18512 12044 18564 12096
rect 19340 12044 19392 12096
rect 19524 12044 19576 12096
rect 23388 12044 23440 12096
rect 29736 12087 29788 12096
rect 29736 12053 29745 12087
rect 29745 12053 29779 12087
rect 29779 12053 29788 12087
rect 29736 12044 29788 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 18144 11840 18196 11892
rect 21456 11840 21508 11892
rect 18052 11772 18104 11824
rect 15568 11747 15620 11756
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 17132 11747 17184 11756
rect 17132 11713 17141 11747
rect 17141 11713 17175 11747
rect 17175 11713 17184 11747
rect 17132 11704 17184 11713
rect 15384 11636 15436 11688
rect 18236 11704 18288 11756
rect 18052 11636 18104 11688
rect 20444 11704 20496 11756
rect 17500 11568 17552 11620
rect 18236 11568 18288 11620
rect 20904 11636 20956 11688
rect 19340 11568 19392 11620
rect 25228 11815 25280 11824
rect 25228 11781 25246 11815
rect 25246 11781 25280 11815
rect 25596 11840 25648 11892
rect 25228 11772 25280 11781
rect 26332 11772 26384 11824
rect 27160 11772 27212 11824
rect 29184 11840 29236 11892
rect 31760 11840 31812 11892
rect 22192 11704 22244 11756
rect 25504 11747 25556 11756
rect 25504 11713 25513 11747
rect 25513 11713 25547 11747
rect 25547 11713 25556 11747
rect 25504 11704 25556 11713
rect 27620 11704 27672 11756
rect 35348 11704 35400 11756
rect 23204 11679 23256 11688
rect 23204 11645 23213 11679
rect 23213 11645 23247 11679
rect 23247 11645 23256 11679
rect 23204 11636 23256 11645
rect 20444 11500 20496 11552
rect 20536 11500 20588 11552
rect 21916 11500 21968 11552
rect 22468 11500 22520 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 14372 11296 14424 11348
rect 13360 11135 13412 11144
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 13360 11092 13412 11101
rect 16212 11296 16264 11348
rect 17592 11296 17644 11348
rect 30380 11339 30432 11348
rect 15384 11160 15436 11212
rect 17868 11228 17920 11280
rect 15200 11092 15252 11144
rect 15936 11135 15988 11144
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 15936 11092 15988 11101
rect 16580 11135 16632 11144
rect 16580 11101 16589 11135
rect 16589 11101 16623 11135
rect 16623 11101 16632 11135
rect 16580 11092 16632 11101
rect 17224 11135 17276 11144
rect 17224 11101 17233 11135
rect 17233 11101 17267 11135
rect 17267 11101 17276 11135
rect 17224 11092 17276 11101
rect 17316 11092 17368 11144
rect 18512 11135 18564 11144
rect 18512 11101 18521 11135
rect 18521 11101 18555 11135
rect 18555 11101 18564 11135
rect 18512 11092 18564 11101
rect 19248 11135 19300 11144
rect 19248 11101 19257 11135
rect 19257 11101 19291 11135
rect 19291 11101 19300 11135
rect 19248 11092 19300 11101
rect 13636 11024 13688 11076
rect 19340 11024 19392 11076
rect 27160 11160 27212 11212
rect 23204 11092 23256 11144
rect 30380 11305 30389 11339
rect 30389 11305 30423 11339
rect 30423 11305 30432 11339
rect 30380 11296 30432 11305
rect 32588 11296 32640 11348
rect 33324 11228 33376 11280
rect 30012 11160 30064 11212
rect 30748 11160 30800 11212
rect 38108 11203 38160 11212
rect 38108 11169 38117 11203
rect 38117 11169 38151 11203
rect 38151 11169 38160 11203
rect 38108 11160 38160 11169
rect 31944 11092 31996 11144
rect 35532 11092 35584 11144
rect 24768 11024 24820 11076
rect 26240 11024 26292 11076
rect 30656 11024 30708 11076
rect 32680 11024 32732 11076
rect 37832 11067 37884 11076
rect 37832 11033 37850 11067
rect 37850 11033 37884 11067
rect 37832 11024 37884 11033
rect 21732 10999 21784 11008
rect 21732 10965 21741 10999
rect 21741 10965 21775 10999
rect 21775 10965 21784 10999
rect 21732 10956 21784 10965
rect 25228 10999 25280 11008
rect 25228 10965 25237 10999
rect 25237 10965 25271 10999
rect 25271 10965 25280 10999
rect 25228 10956 25280 10965
rect 33692 10956 33744 11008
rect 34244 10956 34296 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 15568 10752 15620 10804
rect 19800 10752 19852 10804
rect 19984 10752 20036 10804
rect 15752 10684 15804 10736
rect 21824 10684 21876 10736
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 15476 10659 15528 10668
rect 15476 10625 15485 10659
rect 15485 10625 15519 10659
rect 15519 10625 15528 10659
rect 15476 10616 15528 10625
rect 18328 10616 18380 10668
rect 20076 10659 20128 10668
rect 15384 10548 15436 10600
rect 15568 10548 15620 10600
rect 16856 10548 16908 10600
rect 20076 10625 20085 10659
rect 20085 10625 20119 10659
rect 20119 10625 20128 10659
rect 20076 10616 20128 10625
rect 30196 10752 30248 10804
rect 35532 10727 35584 10736
rect 35532 10693 35541 10727
rect 35541 10693 35575 10727
rect 35575 10693 35584 10727
rect 35532 10684 35584 10693
rect 26056 10616 26108 10668
rect 27160 10616 27212 10668
rect 28356 10616 28408 10668
rect 11704 10523 11756 10532
rect 11704 10489 11713 10523
rect 11713 10489 11747 10523
rect 11747 10489 11756 10523
rect 11704 10480 11756 10489
rect 27620 10548 27672 10600
rect 33784 10659 33836 10668
rect 33784 10625 33793 10659
rect 33793 10625 33827 10659
rect 33827 10625 33836 10659
rect 33784 10616 33836 10625
rect 23204 10480 23256 10532
rect 25504 10480 25556 10532
rect 20260 10455 20312 10464
rect 20260 10421 20269 10455
rect 20269 10421 20303 10455
rect 20303 10421 20312 10455
rect 20260 10412 20312 10421
rect 20444 10412 20496 10464
rect 26424 10412 26476 10464
rect 38016 10455 38068 10464
rect 38016 10421 38025 10455
rect 38025 10421 38059 10455
rect 38059 10421 38068 10455
rect 38016 10412 38068 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 15936 10251 15988 10260
rect 15936 10217 15945 10251
rect 15945 10217 15979 10251
rect 15979 10217 15988 10251
rect 15936 10208 15988 10217
rect 15384 10115 15436 10124
rect 15384 10081 15393 10115
rect 15393 10081 15427 10115
rect 15427 10081 15436 10115
rect 15384 10072 15436 10081
rect 16672 10208 16724 10260
rect 18328 10251 18380 10260
rect 18328 10217 18337 10251
rect 18337 10217 18371 10251
rect 18371 10217 18380 10251
rect 18328 10208 18380 10217
rect 18512 10208 18564 10260
rect 22468 10208 22520 10260
rect 27160 10208 27212 10260
rect 18236 10072 18288 10124
rect 19340 10004 19392 10056
rect 19800 10047 19852 10056
rect 19800 10013 19809 10047
rect 19809 10013 19843 10047
rect 19843 10013 19852 10047
rect 19800 10004 19852 10013
rect 20168 10072 20220 10124
rect 23204 10115 23256 10124
rect 23204 10081 23213 10115
rect 23213 10081 23247 10115
rect 23247 10081 23256 10115
rect 23204 10072 23256 10081
rect 26056 10047 26108 10056
rect 26056 10013 26065 10047
rect 26065 10013 26099 10047
rect 26099 10013 26108 10047
rect 26056 10004 26108 10013
rect 30472 10004 30524 10056
rect 33784 10004 33836 10056
rect 14556 9936 14608 9988
rect 18512 9936 18564 9988
rect 18604 9936 18656 9988
rect 16672 9868 16724 9920
rect 21364 9868 21416 9920
rect 21824 9911 21876 9920
rect 21824 9877 21833 9911
rect 21833 9877 21867 9911
rect 21867 9877 21876 9911
rect 21824 9868 21876 9877
rect 23572 9868 23624 9920
rect 23848 9868 23900 9920
rect 31944 9868 31996 9920
rect 37648 9868 37700 9920
rect 37832 9911 37884 9920
rect 37832 9877 37841 9911
rect 37841 9877 37875 9911
rect 37875 9877 37884 9911
rect 37832 9868 37884 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 11520 9707 11572 9716
rect 11520 9673 11529 9707
rect 11529 9673 11563 9707
rect 11563 9673 11572 9707
rect 11520 9664 11572 9673
rect 18512 9707 18564 9716
rect 18512 9673 18521 9707
rect 18521 9673 18555 9707
rect 18555 9673 18564 9707
rect 18512 9664 18564 9673
rect 9036 9596 9088 9648
rect 10232 9596 10284 9648
rect 11980 9639 12032 9648
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 5816 9528 5868 9580
rect 11980 9460 12032 9512
rect 15292 9596 15344 9648
rect 17776 9596 17828 9648
rect 13452 9528 13504 9580
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 15384 9460 15436 9512
rect 13360 9392 13412 9444
rect 14464 9324 14516 9376
rect 19340 9528 19392 9580
rect 20720 9571 20772 9580
rect 20720 9537 20729 9571
rect 20729 9537 20763 9571
rect 20763 9537 20772 9571
rect 20720 9528 20772 9537
rect 17776 9460 17828 9512
rect 21364 9664 21416 9716
rect 30564 9664 30616 9716
rect 23204 9596 23256 9648
rect 23388 9596 23440 9648
rect 18696 9392 18748 9444
rect 21548 9460 21600 9512
rect 17500 9324 17552 9376
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 22192 9392 22244 9444
rect 25504 9528 25556 9580
rect 23572 9435 23624 9444
rect 23572 9401 23581 9435
rect 23581 9401 23615 9435
rect 23615 9401 23624 9435
rect 23572 9392 23624 9401
rect 24032 9367 24084 9376
rect 24032 9333 24041 9367
rect 24041 9333 24075 9367
rect 24075 9333 24084 9367
rect 24032 9324 24084 9333
rect 24768 9324 24820 9376
rect 28356 9571 28408 9580
rect 28356 9537 28365 9571
rect 28365 9537 28399 9571
rect 28399 9537 28408 9571
rect 28356 9528 28408 9537
rect 26976 9367 27028 9376
rect 26976 9333 26985 9367
rect 26985 9333 27019 9367
rect 27019 9333 27028 9367
rect 26976 9324 27028 9333
rect 27436 9324 27488 9376
rect 31944 9528 31996 9580
rect 35532 9596 35584 9648
rect 34796 9460 34848 9512
rect 29276 9367 29328 9376
rect 29276 9333 29285 9367
rect 29285 9333 29319 9367
rect 29319 9333 29328 9367
rect 29276 9324 29328 9333
rect 29368 9324 29420 9376
rect 35624 9324 35676 9376
rect 37740 9367 37792 9376
rect 37740 9333 37749 9367
rect 37749 9333 37783 9367
rect 37783 9333 37792 9367
rect 37740 9324 37792 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 18604 9120 18656 9172
rect 18696 9163 18748 9172
rect 18696 9129 18705 9163
rect 18705 9129 18739 9163
rect 18739 9129 18748 9163
rect 18696 9120 18748 9129
rect 20720 9120 20772 9172
rect 26424 9163 26476 9172
rect 10416 9052 10468 9104
rect 11980 9052 12032 9104
rect 14832 9095 14884 9104
rect 14832 9061 14841 9095
rect 14841 9061 14875 9095
rect 14875 9061 14884 9095
rect 14832 9052 14884 9061
rect 21548 9052 21600 9104
rect 10232 9027 10284 9036
rect 10232 8993 10241 9027
rect 10241 8993 10275 9027
rect 10275 8993 10284 9027
rect 10232 8984 10284 8993
rect 12440 8984 12492 9036
rect 13912 8916 13964 8968
rect 17500 8959 17552 8968
rect 17500 8925 17509 8959
rect 17509 8925 17543 8959
rect 17543 8925 17552 8959
rect 17500 8916 17552 8925
rect 18696 8984 18748 9036
rect 19340 9027 19392 9036
rect 19340 8993 19349 9027
rect 19349 8993 19383 9027
rect 19383 8993 19392 9027
rect 19340 8984 19392 8993
rect 20536 9027 20588 9036
rect 20536 8993 20545 9027
rect 20545 8993 20579 9027
rect 20579 8993 20588 9027
rect 20536 8984 20588 8993
rect 17868 8916 17920 8968
rect 26424 9129 26433 9163
rect 26433 9129 26467 9163
rect 26467 9129 26476 9163
rect 26424 9120 26476 9129
rect 27344 9120 27396 9172
rect 29184 9120 29236 9172
rect 30656 9120 30708 9172
rect 33232 9163 33284 9172
rect 33232 9129 33241 9163
rect 33241 9129 33275 9163
rect 33275 9129 33284 9163
rect 33232 9120 33284 9129
rect 34796 9120 34848 9172
rect 33600 9052 33652 9104
rect 34336 9052 34388 9104
rect 23204 8984 23256 9036
rect 30564 8916 30616 8968
rect 31944 8959 31996 8968
rect 31944 8925 31953 8959
rect 31953 8925 31987 8959
rect 31987 8925 31996 8959
rect 31944 8916 31996 8925
rect 32404 8916 32456 8968
rect 34704 8959 34756 8968
rect 34704 8925 34713 8959
rect 34713 8925 34747 8959
rect 34747 8925 34756 8959
rect 34704 8916 34756 8925
rect 35532 8916 35584 8968
rect 9864 8848 9916 8900
rect 13268 8848 13320 8900
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 10968 8780 11020 8832
rect 15568 8780 15620 8832
rect 17776 8848 17828 8900
rect 21088 8780 21140 8832
rect 21732 8848 21784 8900
rect 22836 8848 22888 8900
rect 23572 8780 23624 8832
rect 24860 8848 24912 8900
rect 25504 8848 25556 8900
rect 26332 8848 26384 8900
rect 26976 8780 27028 8832
rect 28356 8848 28408 8900
rect 34152 8848 34204 8900
rect 34060 8780 34112 8832
rect 37004 8780 37056 8832
rect 37924 8780 37976 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 12624 8576 12676 8628
rect 13728 8576 13780 8628
rect 13912 8619 13964 8628
rect 13912 8585 13921 8619
rect 13921 8585 13955 8619
rect 13955 8585 13964 8619
rect 13912 8576 13964 8585
rect 14832 8576 14884 8628
rect 15384 8576 15436 8628
rect 15936 8619 15988 8628
rect 15936 8585 15945 8619
rect 15945 8585 15979 8619
rect 15979 8585 15988 8619
rect 15936 8576 15988 8585
rect 16396 8576 16448 8628
rect 20076 8576 20128 8628
rect 8668 8508 8720 8560
rect 10692 8483 10744 8492
rect 10692 8449 10701 8483
rect 10701 8449 10735 8483
rect 10735 8449 10744 8483
rect 10692 8440 10744 8449
rect 11980 8372 12032 8424
rect 14280 8483 14332 8492
rect 14280 8449 14289 8483
rect 14289 8449 14323 8483
rect 14323 8449 14332 8483
rect 14280 8440 14332 8449
rect 16488 8508 16540 8560
rect 17960 8508 18012 8560
rect 20444 8551 20496 8560
rect 15292 8440 15344 8492
rect 15936 8440 15988 8492
rect 20444 8517 20453 8551
rect 20453 8517 20487 8551
rect 20487 8517 20496 8551
rect 20444 8508 20496 8517
rect 22008 8508 22060 8560
rect 29276 8576 29328 8628
rect 34152 8619 34204 8628
rect 34152 8585 34161 8619
rect 34161 8585 34195 8619
rect 34195 8585 34204 8619
rect 34152 8576 34204 8585
rect 35440 8576 35492 8628
rect 34612 8508 34664 8560
rect 35808 8551 35860 8560
rect 35808 8517 35817 8551
rect 35817 8517 35851 8551
rect 35851 8517 35860 8551
rect 35808 8508 35860 8517
rect 17684 8372 17736 8424
rect 19984 8372 20036 8424
rect 20076 8372 20128 8424
rect 20444 8372 20496 8424
rect 21088 8372 21140 8424
rect 21272 8372 21324 8424
rect 22376 8440 22428 8492
rect 23204 8483 23256 8492
rect 23204 8449 23213 8483
rect 23213 8449 23247 8483
rect 23247 8449 23256 8483
rect 23204 8440 23256 8449
rect 26240 8440 26292 8492
rect 28356 8483 28408 8492
rect 28356 8449 28365 8483
rect 28365 8449 28399 8483
rect 28399 8449 28408 8483
rect 28356 8440 28408 8449
rect 34428 8440 34480 8492
rect 21732 8304 21784 8356
rect 15384 8236 15436 8288
rect 20444 8236 20496 8288
rect 26148 8304 26200 8356
rect 22008 8236 22060 8288
rect 27436 8236 27488 8288
rect 30656 8304 30708 8356
rect 37372 8347 37424 8356
rect 37372 8313 37381 8347
rect 37381 8313 37415 8347
rect 37415 8313 37424 8347
rect 37372 8304 37424 8313
rect 38108 8304 38160 8356
rect 32220 8279 32272 8288
rect 32220 8245 32229 8279
rect 32229 8245 32263 8279
rect 32263 8245 32272 8279
rect 32220 8236 32272 8245
rect 35348 8236 35400 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 10324 8032 10376 8084
rect 12624 8075 12676 8084
rect 12624 8041 12633 8075
rect 12633 8041 12667 8075
rect 12667 8041 12676 8075
rect 12624 8032 12676 8041
rect 24860 8032 24912 8084
rect 30472 8075 30524 8084
rect 30472 8041 30481 8075
rect 30481 8041 30515 8075
rect 30515 8041 30524 8075
rect 30472 8032 30524 8041
rect 30840 8032 30892 8084
rect 33968 8032 34020 8084
rect 34704 8075 34756 8084
rect 34704 8041 34713 8075
rect 34713 8041 34747 8075
rect 34747 8041 34756 8075
rect 34704 8032 34756 8041
rect 37096 8032 37148 8084
rect 15108 7964 15160 8016
rect 11152 7896 11204 7948
rect 15200 7871 15252 7880
rect 15200 7837 15209 7871
rect 15209 7837 15243 7871
rect 15243 7837 15252 7871
rect 15200 7828 15252 7837
rect 15384 7871 15436 7880
rect 15384 7837 15393 7871
rect 15393 7837 15427 7871
rect 15427 7837 15436 7871
rect 15384 7828 15436 7837
rect 17960 7896 18012 7948
rect 19340 7896 19392 7948
rect 20444 7896 20496 7948
rect 17408 7828 17460 7880
rect 18696 7828 18748 7880
rect 19248 7871 19300 7880
rect 19248 7837 19257 7871
rect 19257 7837 19291 7871
rect 19291 7837 19300 7871
rect 19248 7828 19300 7837
rect 32404 7939 32456 7948
rect 32404 7905 32413 7939
rect 32413 7905 32447 7939
rect 32447 7905 32456 7939
rect 32404 7896 32456 7905
rect 35624 7964 35676 8016
rect 35348 7939 35400 7948
rect 35348 7905 35357 7939
rect 35357 7905 35391 7939
rect 35391 7905 35400 7939
rect 35348 7896 35400 7905
rect 12072 7760 12124 7812
rect 19340 7760 19392 7812
rect 17040 7692 17092 7744
rect 20812 7692 20864 7744
rect 22284 7760 22336 7812
rect 23480 7828 23532 7880
rect 27620 7871 27672 7880
rect 27620 7837 27629 7871
rect 27629 7837 27663 7871
rect 27663 7837 27672 7871
rect 27620 7828 27672 7837
rect 32220 7828 32272 7880
rect 29092 7760 29144 7812
rect 34796 7828 34848 7880
rect 36176 7828 36228 7880
rect 38200 7828 38252 7880
rect 23756 7692 23808 7744
rect 26240 7735 26292 7744
rect 26240 7701 26249 7735
rect 26249 7701 26283 7735
rect 26283 7701 26292 7735
rect 26240 7692 26292 7701
rect 33140 7692 33192 7744
rect 35808 7692 35860 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 10324 7488 10376 7540
rect 12072 7531 12124 7540
rect 12072 7497 12081 7531
rect 12081 7497 12115 7531
rect 12115 7497 12124 7531
rect 12072 7488 12124 7497
rect 15200 7488 15252 7540
rect 15936 7488 15988 7540
rect 16948 7531 17000 7540
rect 16948 7497 16957 7531
rect 16957 7497 16991 7531
rect 16991 7497 17000 7531
rect 16948 7488 17000 7497
rect 17408 7531 17460 7540
rect 17408 7497 17417 7531
rect 17417 7497 17451 7531
rect 17451 7497 17460 7531
rect 17408 7488 17460 7497
rect 18696 7531 18748 7540
rect 18696 7497 18705 7531
rect 18705 7497 18739 7531
rect 18739 7497 18748 7531
rect 18696 7488 18748 7497
rect 7012 7420 7064 7472
rect 9956 7352 10008 7404
rect 12164 7352 12216 7404
rect 13544 7395 13596 7404
rect 13544 7361 13553 7395
rect 13553 7361 13587 7395
rect 13587 7361 13596 7395
rect 13544 7352 13596 7361
rect 13728 7395 13780 7404
rect 13728 7361 13737 7395
rect 13737 7361 13771 7395
rect 13771 7361 13780 7395
rect 13728 7352 13780 7361
rect 15292 7420 15344 7472
rect 20720 7488 20772 7540
rect 26240 7488 26292 7540
rect 29092 7531 29144 7540
rect 29092 7497 29101 7531
rect 29101 7497 29135 7531
rect 29135 7497 29144 7531
rect 29092 7488 29144 7497
rect 34796 7531 34848 7540
rect 10416 7327 10468 7336
rect 10416 7293 10425 7327
rect 10425 7293 10459 7327
rect 10459 7293 10468 7327
rect 10416 7284 10468 7293
rect 12624 7284 12676 7336
rect 14464 7284 14516 7336
rect 15476 7352 15528 7404
rect 18512 7352 18564 7404
rect 15936 7284 15988 7336
rect 16488 7284 16540 7336
rect 18144 7327 18196 7336
rect 18144 7293 18153 7327
rect 18153 7293 18187 7327
rect 18187 7293 18196 7327
rect 18144 7284 18196 7293
rect 34796 7497 34805 7531
rect 34805 7497 34839 7531
rect 34839 7497 34848 7531
rect 34796 7488 34848 7497
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 30380 7420 30432 7472
rect 37096 7488 37148 7540
rect 37280 7420 37332 7472
rect 30288 7352 30340 7404
rect 32128 7395 32180 7404
rect 32128 7361 32137 7395
rect 32137 7361 32171 7395
rect 32171 7361 32180 7395
rect 32128 7352 32180 7361
rect 33416 7352 33468 7404
rect 33968 7352 34020 7404
rect 17960 7216 18012 7268
rect 23480 7284 23532 7336
rect 31484 7284 31536 7336
rect 20720 7216 20772 7268
rect 11520 7148 11572 7200
rect 12624 7148 12676 7200
rect 14096 7148 14148 7200
rect 17500 7148 17552 7200
rect 31300 7148 31352 7200
rect 32312 7191 32364 7200
rect 32312 7157 32321 7191
rect 32321 7157 32355 7191
rect 32355 7157 32364 7191
rect 32312 7148 32364 7157
rect 32772 7191 32824 7200
rect 32772 7157 32781 7191
rect 32781 7157 32815 7191
rect 32815 7157 32824 7191
rect 32772 7148 32824 7157
rect 35992 7352 36044 7404
rect 34060 7216 34112 7268
rect 35900 7216 35952 7268
rect 35348 7148 35400 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 15936 6987 15988 6996
rect 15936 6953 15945 6987
rect 15945 6953 15979 6987
rect 15979 6953 15988 6987
rect 15936 6944 15988 6953
rect 12440 6808 12492 6860
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 12348 6740 12400 6792
rect 12624 6672 12676 6724
rect 14096 6808 14148 6860
rect 14464 6851 14516 6860
rect 14464 6817 14473 6851
rect 14473 6817 14507 6851
rect 14507 6817 14516 6851
rect 14464 6808 14516 6817
rect 15568 6808 15620 6860
rect 16948 6944 17000 6996
rect 19248 6987 19300 6996
rect 19248 6953 19257 6987
rect 19257 6953 19291 6987
rect 19291 6953 19300 6987
rect 19248 6944 19300 6953
rect 19340 6876 19392 6928
rect 19156 6808 19208 6860
rect 21732 6808 21784 6860
rect 30564 6851 30616 6860
rect 13912 6740 13964 6792
rect 20076 6740 20128 6792
rect 22192 6740 22244 6792
rect 16396 6672 16448 6724
rect 19340 6672 19392 6724
rect 19524 6672 19576 6724
rect 11060 6647 11112 6656
rect 11060 6613 11069 6647
rect 11069 6613 11103 6647
rect 11103 6613 11112 6647
rect 11060 6604 11112 6613
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 17408 6647 17460 6656
rect 17408 6613 17417 6647
rect 17417 6613 17451 6647
rect 17451 6613 17460 6647
rect 17408 6604 17460 6613
rect 18972 6604 19024 6656
rect 20168 6604 20220 6656
rect 22284 6672 22336 6724
rect 21640 6647 21692 6656
rect 21640 6613 21649 6647
rect 21649 6613 21683 6647
rect 21683 6613 21692 6647
rect 21640 6604 21692 6613
rect 21732 6604 21784 6656
rect 23480 6740 23532 6792
rect 23572 6740 23624 6792
rect 27620 6740 27672 6792
rect 28356 6740 28408 6792
rect 24768 6672 24820 6724
rect 30564 6817 30573 6851
rect 30573 6817 30607 6851
rect 30607 6817 30616 6851
rect 30564 6808 30616 6817
rect 30748 6851 30800 6860
rect 30748 6817 30757 6851
rect 30757 6817 30791 6851
rect 30791 6817 30800 6851
rect 30748 6808 30800 6817
rect 34336 6808 34388 6860
rect 35348 6851 35400 6860
rect 35348 6817 35357 6851
rect 35357 6817 35391 6851
rect 35391 6817 35400 6851
rect 35348 6808 35400 6817
rect 36176 6851 36228 6860
rect 36176 6817 36185 6851
rect 36185 6817 36219 6851
rect 36219 6817 36228 6851
rect 36176 6808 36228 6817
rect 31484 6740 31536 6792
rect 33968 6783 34020 6792
rect 33968 6749 33977 6783
rect 33977 6749 34011 6783
rect 34011 6749 34020 6783
rect 33968 6740 34020 6749
rect 37188 6740 37240 6792
rect 30840 6647 30892 6656
rect 30840 6613 30849 6647
rect 30849 6613 30883 6647
rect 30883 6613 30892 6647
rect 30840 6604 30892 6613
rect 32312 6672 32364 6724
rect 32128 6604 32180 6656
rect 34428 6604 34480 6656
rect 36084 6604 36136 6656
rect 37556 6647 37608 6656
rect 37556 6613 37565 6647
rect 37565 6613 37599 6647
rect 37599 6613 37608 6647
rect 37556 6604 37608 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 9680 6400 9732 6452
rect 8392 6332 8444 6384
rect 12164 6400 12216 6452
rect 13912 6443 13964 6452
rect 13912 6409 13921 6443
rect 13921 6409 13955 6443
rect 13955 6409 13964 6443
rect 13912 6400 13964 6409
rect 18972 6443 19024 6452
rect 10416 6332 10468 6384
rect 12072 6332 12124 6384
rect 12532 6332 12584 6384
rect 13360 6332 13412 6384
rect 11704 6264 11756 6316
rect 12624 6264 12676 6316
rect 12900 6307 12952 6316
rect 12900 6273 12909 6307
rect 12909 6273 12943 6307
rect 12943 6273 12952 6307
rect 12900 6264 12952 6273
rect 13176 6264 13228 6316
rect 13544 6307 13596 6316
rect 13544 6273 13553 6307
rect 13553 6273 13587 6307
rect 13587 6273 13596 6307
rect 13544 6264 13596 6273
rect 12348 6196 12400 6248
rect 13728 6307 13780 6316
rect 13728 6273 13737 6307
rect 13737 6273 13771 6307
rect 13771 6273 13780 6307
rect 16488 6332 16540 6384
rect 13728 6264 13780 6273
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 18972 6409 18981 6443
rect 18981 6409 19015 6443
rect 19015 6409 19024 6443
rect 18972 6400 19024 6409
rect 19340 6400 19392 6452
rect 20168 6443 20220 6452
rect 20168 6409 20177 6443
rect 20177 6409 20211 6443
rect 20211 6409 20220 6443
rect 20168 6400 20220 6409
rect 22284 6400 22336 6452
rect 22376 6400 22428 6452
rect 28816 6400 28868 6452
rect 30288 6443 30340 6452
rect 18144 6332 18196 6384
rect 28356 6332 28408 6384
rect 30288 6409 30297 6443
rect 30297 6409 30331 6443
rect 30331 6409 30340 6443
rect 30288 6400 30340 6409
rect 31392 6400 31444 6452
rect 32496 6400 32548 6452
rect 33968 6400 34020 6452
rect 34336 6400 34388 6452
rect 16120 6264 16172 6273
rect 17040 6264 17092 6316
rect 16856 6196 16908 6248
rect 17776 6196 17828 6248
rect 17316 6128 17368 6180
rect 18604 6264 18656 6316
rect 29000 6264 29052 6316
rect 30564 6332 30616 6384
rect 30656 6307 30708 6316
rect 30656 6273 30665 6307
rect 30665 6273 30699 6307
rect 30699 6273 30708 6307
rect 30656 6264 30708 6273
rect 23480 6196 23532 6248
rect 32036 6196 32088 6248
rect 33232 6332 33284 6384
rect 33968 6264 34020 6316
rect 34704 6264 34756 6316
rect 33692 6196 33744 6248
rect 12532 6060 12584 6112
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 15752 6103 15804 6112
rect 15752 6069 15761 6103
rect 15761 6069 15795 6103
rect 15795 6069 15804 6103
rect 15752 6060 15804 6069
rect 16396 6060 16448 6112
rect 20260 6128 20312 6180
rect 20444 6128 20496 6180
rect 21456 6128 21508 6180
rect 17776 6060 17828 6112
rect 21824 6103 21876 6112
rect 21824 6069 21833 6103
rect 21833 6069 21867 6103
rect 21867 6069 21876 6103
rect 21824 6060 21876 6069
rect 32956 6128 33008 6180
rect 24768 6060 24820 6112
rect 24860 6060 24912 6112
rect 32496 6060 32548 6112
rect 37556 6128 37608 6180
rect 34796 6103 34848 6112
rect 34796 6069 34805 6103
rect 34805 6069 34839 6103
rect 34839 6069 34848 6103
rect 34796 6060 34848 6069
rect 35348 6103 35400 6112
rect 35348 6069 35357 6103
rect 35357 6069 35391 6103
rect 35391 6069 35400 6103
rect 35348 6060 35400 6069
rect 36636 6060 36688 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 9956 5899 10008 5908
rect 9956 5865 9965 5899
rect 9965 5865 9999 5899
rect 9999 5865 10008 5899
rect 9956 5856 10008 5865
rect 12072 5899 12124 5908
rect 12072 5865 12081 5899
rect 12081 5865 12115 5899
rect 12115 5865 12124 5899
rect 12072 5856 12124 5865
rect 12900 5899 12952 5908
rect 12900 5865 12909 5899
rect 12909 5865 12943 5899
rect 12943 5865 12952 5899
rect 12900 5856 12952 5865
rect 12992 5856 13044 5908
rect 16120 5856 16172 5908
rect 19432 5856 19484 5908
rect 18604 5788 18656 5840
rect 19340 5788 19392 5840
rect 20536 5831 20588 5840
rect 20536 5797 20545 5831
rect 20545 5797 20579 5831
rect 20579 5797 20588 5831
rect 20536 5788 20588 5797
rect 9680 5720 9732 5772
rect 13176 5720 13228 5772
rect 15752 5720 15804 5772
rect 16488 5720 16540 5772
rect 17500 5720 17552 5772
rect 10416 5652 10468 5704
rect 10876 5695 10928 5704
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 12716 5652 12768 5704
rect 14096 5652 14148 5704
rect 16856 5652 16908 5704
rect 17316 5652 17368 5704
rect 26148 5856 26200 5908
rect 31392 5899 31444 5908
rect 31392 5865 31401 5899
rect 31401 5865 31435 5899
rect 31435 5865 31444 5899
rect 31392 5856 31444 5865
rect 33140 5856 33192 5908
rect 33232 5856 33284 5908
rect 34704 5899 34756 5908
rect 34704 5865 34713 5899
rect 34713 5865 34747 5899
rect 34747 5865 34756 5899
rect 34704 5856 34756 5865
rect 35992 5899 36044 5908
rect 35992 5865 36001 5899
rect 36001 5865 36035 5899
rect 36035 5865 36044 5899
rect 35992 5856 36044 5865
rect 29184 5788 29236 5840
rect 32036 5831 32088 5840
rect 32036 5797 32045 5831
rect 32045 5797 32079 5831
rect 32079 5797 32088 5831
rect 32036 5788 32088 5797
rect 37372 5856 37424 5908
rect 36176 5788 36228 5840
rect 35348 5763 35400 5772
rect 35348 5729 35357 5763
rect 35357 5729 35391 5763
rect 35391 5729 35400 5763
rect 35348 5720 35400 5729
rect 21272 5695 21324 5704
rect 21272 5661 21281 5695
rect 21281 5661 21315 5695
rect 21315 5661 21324 5695
rect 21272 5652 21324 5661
rect 21456 5695 21508 5704
rect 21456 5661 21465 5695
rect 21465 5661 21499 5695
rect 21499 5661 21508 5695
rect 21456 5652 21508 5661
rect 22652 5652 22704 5704
rect 23480 5695 23532 5704
rect 23480 5661 23489 5695
rect 23489 5661 23523 5695
rect 23523 5661 23532 5695
rect 23480 5652 23532 5661
rect 27620 5652 27672 5704
rect 28356 5652 28408 5704
rect 29644 5652 29696 5704
rect 8484 5584 8536 5636
rect 14004 5584 14056 5636
rect 14464 5584 14516 5636
rect 8300 5516 8352 5568
rect 12532 5516 12584 5568
rect 14740 5516 14792 5568
rect 17500 5584 17552 5636
rect 17960 5627 18012 5636
rect 17960 5593 17969 5627
rect 17969 5593 18003 5627
rect 18003 5593 18012 5627
rect 17960 5584 18012 5593
rect 18236 5584 18288 5636
rect 19340 5584 19392 5636
rect 20260 5584 20312 5636
rect 22284 5584 22336 5636
rect 23664 5584 23716 5636
rect 25044 5584 25096 5636
rect 27344 5584 27396 5636
rect 29184 5584 29236 5636
rect 31484 5652 31536 5704
rect 35900 5652 35952 5704
rect 32588 5584 32640 5636
rect 34796 5584 34848 5636
rect 17224 5516 17276 5568
rect 19432 5516 19484 5568
rect 20720 5559 20772 5568
rect 20720 5525 20729 5559
rect 20729 5525 20763 5559
rect 20763 5525 20772 5559
rect 20720 5516 20772 5525
rect 32496 5559 32548 5568
rect 32496 5525 32505 5559
rect 32505 5525 32539 5559
rect 32539 5525 32548 5559
rect 32496 5516 32548 5525
rect 34520 5516 34572 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 10508 5355 10560 5364
rect 10508 5321 10517 5355
rect 10517 5321 10551 5355
rect 10551 5321 10560 5355
rect 10508 5312 10560 5321
rect 10876 5312 10928 5364
rect 10324 5244 10376 5296
rect 15016 5312 15068 5364
rect 15568 5312 15620 5364
rect 19064 5355 19116 5364
rect 19064 5321 19073 5355
rect 19073 5321 19107 5355
rect 19107 5321 19116 5355
rect 19064 5312 19116 5321
rect 19984 5312 20036 5364
rect 20720 5312 20772 5364
rect 9680 5176 9732 5228
rect 10968 5176 11020 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 12164 5176 12216 5228
rect 13820 5244 13872 5296
rect 17224 5244 17276 5296
rect 21272 5244 21324 5296
rect 21916 5244 21968 5296
rect 24952 5244 25004 5296
rect 25596 5287 25648 5296
rect 25596 5253 25605 5287
rect 25605 5253 25639 5287
rect 25639 5253 25648 5287
rect 25596 5244 25648 5253
rect 26332 5244 26384 5296
rect 26516 5244 26568 5296
rect 27712 5244 27764 5296
rect 15568 5219 15620 5228
rect 10048 5108 10100 5160
rect 10416 5151 10468 5160
rect 10416 5117 10425 5151
rect 10425 5117 10459 5151
rect 10459 5117 10468 5151
rect 10416 5108 10468 5117
rect 12808 5108 12860 5160
rect 13544 5108 13596 5160
rect 14924 5151 14976 5160
rect 14924 5117 14933 5151
rect 14933 5117 14967 5151
rect 14967 5117 14976 5151
rect 14924 5108 14976 5117
rect 15568 5185 15577 5219
rect 15577 5185 15611 5219
rect 15611 5185 15620 5219
rect 15568 5176 15620 5185
rect 15660 5176 15712 5228
rect 16396 5176 16448 5228
rect 16488 5108 16540 5160
rect 17040 5151 17092 5160
rect 17040 5117 17049 5151
rect 17049 5117 17083 5151
rect 17083 5117 17092 5151
rect 17040 5108 17092 5117
rect 17408 5176 17460 5228
rect 18880 5219 18932 5228
rect 18880 5185 18889 5219
rect 18889 5185 18923 5219
rect 18923 5185 18932 5219
rect 18880 5176 18932 5185
rect 19340 5176 19392 5228
rect 24860 5176 24912 5228
rect 27804 5176 27856 5228
rect 7840 5040 7892 5092
rect 10692 5040 10744 5092
rect 17960 5108 18012 5160
rect 23480 5151 23532 5160
rect 17316 5040 17368 5092
rect 18328 5040 18380 5092
rect 23480 5117 23489 5151
rect 23489 5117 23523 5151
rect 23523 5117 23532 5151
rect 23480 5108 23532 5117
rect 28356 5151 28408 5160
rect 28356 5117 28365 5151
rect 28365 5117 28399 5151
rect 28399 5117 28408 5151
rect 28356 5108 28408 5117
rect 32496 5108 32548 5160
rect 33600 5244 33652 5296
rect 33784 5287 33836 5296
rect 33784 5253 33793 5287
rect 33793 5253 33827 5287
rect 33827 5253 33836 5287
rect 33784 5244 33836 5253
rect 36176 5244 36228 5296
rect 36912 5312 36964 5364
rect 37372 5244 37424 5296
rect 7564 5015 7616 5024
rect 7564 4981 7573 5015
rect 7573 4981 7607 5015
rect 7607 4981 7616 5015
rect 7564 4972 7616 4981
rect 10508 4972 10560 5024
rect 10968 4972 11020 5024
rect 12164 4972 12216 5024
rect 13084 5015 13136 5024
rect 13084 4981 13093 5015
rect 13093 4981 13127 5015
rect 13127 4981 13136 5015
rect 13084 4972 13136 4981
rect 14188 4972 14240 5024
rect 14372 4972 14424 5024
rect 15108 5015 15160 5024
rect 15108 4981 15117 5015
rect 15117 4981 15151 5015
rect 15151 4981 15160 5015
rect 15108 4972 15160 4981
rect 15844 5015 15896 5024
rect 15844 4981 15853 5015
rect 15853 4981 15887 5015
rect 15887 4981 15896 5015
rect 15844 4972 15896 4981
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 21824 5015 21876 5024
rect 21824 4981 21833 5015
rect 21833 4981 21867 5015
rect 21867 4981 21876 5015
rect 21824 4972 21876 4981
rect 28724 4972 28776 5024
rect 29736 5040 29788 5092
rect 32864 5108 32916 5160
rect 33048 5040 33100 5092
rect 37464 5219 37516 5228
rect 37464 5185 37473 5219
rect 37473 5185 37507 5219
rect 37507 5185 37516 5219
rect 37464 5176 37516 5185
rect 38108 5219 38160 5228
rect 38108 5185 38117 5219
rect 38117 5185 38151 5219
rect 38151 5185 38160 5219
rect 38108 5176 38160 5185
rect 36452 5040 36504 5092
rect 29368 5015 29420 5024
rect 29368 4981 29377 5015
rect 29377 4981 29411 5015
rect 29411 4981 29420 5015
rect 29368 4972 29420 4981
rect 29828 4972 29880 5024
rect 30564 5015 30616 5024
rect 30564 4981 30573 5015
rect 30573 4981 30607 5015
rect 30607 4981 30616 5015
rect 30564 4972 30616 4981
rect 31576 5015 31628 5024
rect 31576 4981 31585 5015
rect 31585 4981 31619 5015
rect 31619 4981 31628 5015
rect 31576 4972 31628 4981
rect 36268 4972 36320 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 12624 4768 12676 4820
rect 9404 4743 9456 4752
rect 9404 4709 9413 4743
rect 9413 4709 9447 4743
rect 9447 4709 9456 4743
rect 9404 4700 9456 4709
rect 10140 4632 10192 4684
rect 13728 4700 13780 4752
rect 15568 4768 15620 4820
rect 16488 4811 16540 4820
rect 16488 4777 16497 4811
rect 16497 4777 16531 4811
rect 16531 4777 16540 4811
rect 16488 4768 16540 4777
rect 16948 4768 17000 4820
rect 17500 4768 17552 4820
rect 19432 4768 19484 4820
rect 20168 4768 20220 4820
rect 20260 4768 20312 4820
rect 21088 4768 21140 4820
rect 21272 4768 21324 4820
rect 14924 4700 14976 4752
rect 17040 4700 17092 4752
rect 24584 4768 24636 4820
rect 33692 4768 33744 4820
rect 34520 4768 34572 4820
rect 37464 4768 37516 4820
rect 9496 4564 9548 4616
rect 10416 4607 10468 4616
rect 10416 4573 10425 4607
rect 10425 4573 10459 4607
rect 10459 4573 10468 4607
rect 10416 4564 10468 4573
rect 12716 4607 12768 4616
rect 12716 4573 12725 4607
rect 12725 4573 12759 4607
rect 12759 4573 12768 4607
rect 12716 4564 12768 4573
rect 12992 4564 13044 4616
rect 13268 4564 13320 4616
rect 14188 4607 14240 4616
rect 14188 4573 14197 4607
rect 14197 4573 14231 4607
rect 14231 4573 14240 4607
rect 14188 4564 14240 4573
rect 14372 4607 14424 4616
rect 14372 4573 14381 4607
rect 14381 4573 14415 4607
rect 14415 4573 14424 4607
rect 14372 4564 14424 4573
rect 15108 4632 15160 4684
rect 18604 4632 18656 4684
rect 32036 4700 32088 4752
rect 15660 4564 15712 4616
rect 18052 4564 18104 4616
rect 8116 4496 8168 4548
rect 5264 4471 5316 4480
rect 5264 4437 5273 4471
rect 5273 4437 5307 4471
rect 5307 4437 5316 4471
rect 5264 4428 5316 4437
rect 5632 4428 5684 4480
rect 10968 4428 11020 4480
rect 11980 4428 12032 4480
rect 12256 4471 12308 4480
rect 12256 4437 12265 4471
rect 12265 4437 12299 4471
rect 12299 4437 12308 4471
rect 12256 4428 12308 4437
rect 15936 4496 15988 4548
rect 19432 4564 19484 4616
rect 20536 4564 20588 4616
rect 23480 4564 23532 4616
rect 23572 4564 23624 4616
rect 31576 4632 31628 4684
rect 27068 4564 27120 4616
rect 28356 4564 28408 4616
rect 32128 4564 32180 4616
rect 33048 4632 33100 4684
rect 35348 4700 35400 4752
rect 37372 4743 37424 4752
rect 37372 4709 37381 4743
rect 37381 4709 37415 4743
rect 37415 4709 37424 4743
rect 37372 4700 37424 4709
rect 35440 4632 35492 4684
rect 32680 4564 32732 4616
rect 32956 4607 33008 4616
rect 32956 4573 32965 4607
rect 32965 4573 32999 4607
rect 32999 4573 33008 4607
rect 32956 4564 33008 4573
rect 33876 4564 33928 4616
rect 34060 4564 34112 4616
rect 36084 4564 36136 4616
rect 36268 4607 36320 4616
rect 36268 4573 36302 4607
rect 36302 4573 36320 4607
rect 36268 4564 36320 4573
rect 37924 4564 37976 4616
rect 15200 4428 15252 4480
rect 16856 4428 16908 4480
rect 19248 4428 19300 4480
rect 20444 4428 20496 4480
rect 21272 4428 21324 4480
rect 21640 4471 21692 4480
rect 21640 4437 21649 4471
rect 21649 4437 21683 4471
rect 21683 4437 21692 4471
rect 21640 4428 21692 4437
rect 22376 4496 22428 4548
rect 23848 4496 23900 4548
rect 26424 4496 26476 4548
rect 31208 4496 31260 4548
rect 22100 4428 22152 4480
rect 27160 4428 27212 4480
rect 29000 4471 29052 4480
rect 29000 4437 29009 4471
rect 29009 4437 29043 4471
rect 29043 4437 29052 4471
rect 29000 4428 29052 4437
rect 29920 4471 29972 4480
rect 29920 4437 29929 4471
rect 29929 4437 29963 4471
rect 29963 4437 29972 4471
rect 29920 4428 29972 4437
rect 36544 4496 36596 4548
rect 33140 4471 33192 4480
rect 33140 4437 33149 4471
rect 33149 4437 33183 4471
rect 33183 4437 33192 4471
rect 33140 4428 33192 4437
rect 35072 4471 35124 4480
rect 35072 4437 35081 4471
rect 35081 4437 35115 4471
rect 35115 4437 35124 4471
rect 35072 4428 35124 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 8576 4224 8628 4276
rect 9404 4224 9456 4276
rect 10416 4224 10468 4276
rect 10692 4224 10744 4276
rect 12992 4224 13044 4276
rect 15660 4224 15712 4276
rect 17776 4224 17828 4276
rect 18420 4224 18472 4276
rect 23572 4224 23624 4276
rect 28448 4267 28500 4276
rect 28448 4233 28457 4267
rect 28457 4233 28491 4267
rect 28491 4233 28500 4267
rect 28448 4224 28500 4233
rect 10232 4131 10284 4140
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10232 4088 10284 4097
rect 11520 4088 11572 4140
rect 12072 4131 12124 4140
rect 12072 4097 12081 4131
rect 12081 4097 12115 4131
rect 12115 4097 12124 4131
rect 12072 4088 12124 4097
rect 12440 4088 12492 4140
rect 12900 4156 12952 4208
rect 12716 4131 12768 4140
rect 12716 4097 12725 4131
rect 12725 4097 12759 4131
rect 12759 4097 12768 4131
rect 12716 4088 12768 4097
rect 9036 4020 9088 4072
rect 10048 4063 10100 4072
rect 10048 4029 10057 4063
rect 10057 4029 10091 4063
rect 10091 4029 10100 4063
rect 10048 4020 10100 4029
rect 10416 4020 10468 4072
rect 13544 4131 13596 4140
rect 13544 4097 13553 4131
rect 13553 4097 13587 4131
rect 13587 4097 13596 4131
rect 13544 4088 13596 4097
rect 13728 4088 13780 4140
rect 13820 4020 13872 4072
rect 16488 4156 16540 4208
rect 14740 4088 14792 4140
rect 15568 4088 15620 4140
rect 16856 4088 16908 4140
rect 17224 4131 17276 4140
rect 17224 4097 17233 4131
rect 17233 4097 17267 4131
rect 17267 4097 17276 4131
rect 17224 4088 17276 4097
rect 17592 4131 17644 4140
rect 17592 4097 17601 4131
rect 17601 4097 17635 4131
rect 17635 4097 17644 4131
rect 17592 4088 17644 4097
rect 17776 4131 17828 4140
rect 17776 4097 17785 4131
rect 17785 4097 17819 4131
rect 17819 4097 17828 4131
rect 17776 4088 17828 4097
rect 15844 4020 15896 4072
rect 16396 4020 16448 4072
rect 17960 4020 18012 4072
rect 7288 3952 7340 4004
rect 10600 3952 10652 4004
rect 4068 3884 4120 3936
rect 4620 3927 4672 3936
rect 4620 3893 4629 3927
rect 4629 3893 4663 3927
rect 4663 3893 4672 3927
rect 4620 3884 4672 3893
rect 5540 3884 5592 3936
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 9404 3927 9456 3936
rect 9404 3893 9413 3927
rect 9413 3893 9447 3927
rect 9447 3893 9456 3927
rect 9404 3884 9456 3893
rect 9588 3884 9640 3936
rect 12440 3952 12492 4004
rect 12808 3952 12860 4004
rect 12256 3927 12308 3936
rect 12256 3893 12265 3927
rect 12265 3893 12299 3927
rect 12299 3893 12308 3927
rect 12256 3884 12308 3893
rect 14280 3952 14332 4004
rect 15752 3952 15804 4004
rect 18328 4088 18380 4140
rect 19340 4088 19392 4140
rect 21088 4156 21140 4208
rect 23940 4156 23992 4208
rect 31208 4224 31260 4276
rect 31668 4224 31720 4276
rect 32128 4267 32180 4276
rect 32128 4233 32137 4267
rect 32137 4233 32171 4267
rect 32171 4233 32180 4267
rect 32128 4224 32180 4233
rect 33140 4224 33192 4276
rect 35072 4224 35124 4276
rect 35440 4224 35492 4276
rect 29920 4156 29972 4208
rect 32496 4199 32548 4208
rect 32496 4165 32505 4199
rect 32505 4165 32539 4199
rect 32539 4165 32548 4199
rect 32496 4156 32548 4165
rect 33048 4156 33100 4208
rect 19984 4088 20036 4140
rect 21180 4131 21232 4140
rect 21180 4097 21189 4131
rect 21189 4097 21223 4131
rect 21223 4097 21232 4131
rect 21180 4088 21232 4097
rect 21272 4088 21324 4140
rect 22744 4088 22796 4140
rect 23480 4088 23532 4140
rect 24216 4088 24268 4140
rect 27160 4088 27212 4140
rect 28264 4088 28316 4140
rect 29000 4088 29052 4140
rect 32588 4131 32640 4140
rect 24032 4020 24084 4072
rect 27068 4063 27120 4072
rect 27068 4029 27077 4063
rect 27077 4029 27111 4063
rect 27111 4029 27120 4063
rect 27068 4020 27120 4029
rect 28448 4020 28500 4072
rect 20076 3995 20128 4004
rect 20076 3961 20085 3995
rect 20085 3961 20119 3995
rect 20119 3961 20128 3995
rect 20076 3952 20128 3961
rect 20168 3952 20220 4004
rect 21824 3995 21876 4004
rect 21824 3961 21833 3995
rect 21833 3961 21867 3995
rect 21867 3961 21876 3995
rect 21824 3952 21876 3961
rect 14372 3884 14424 3936
rect 15476 3884 15528 3936
rect 15844 3927 15896 3936
rect 15844 3893 15853 3927
rect 15853 3893 15887 3927
rect 15887 3893 15896 3927
rect 15844 3884 15896 3893
rect 16764 3927 16816 3936
rect 16764 3893 16773 3927
rect 16773 3893 16807 3927
rect 16807 3893 16816 3927
rect 16764 3884 16816 3893
rect 21088 3884 21140 3936
rect 21272 3884 21324 3936
rect 26240 3952 26292 4004
rect 26976 3952 27028 4004
rect 32588 4097 32597 4131
rect 32597 4097 32631 4131
rect 32631 4097 32640 4131
rect 32588 4088 32640 4097
rect 32036 4020 32088 4072
rect 33048 4020 33100 4072
rect 36084 4156 36136 4208
rect 36360 4156 36412 4208
rect 33232 4088 33284 4140
rect 35992 4088 36044 4140
rect 36452 4131 36504 4140
rect 36452 4097 36470 4131
rect 36470 4097 36504 4131
rect 36452 4088 36504 4097
rect 35716 4020 35768 4072
rect 22468 3927 22520 3936
rect 22468 3893 22477 3927
rect 22477 3893 22511 3927
rect 22511 3893 22520 3927
rect 22468 3884 22520 3893
rect 22836 3884 22888 3936
rect 23204 3884 23256 3936
rect 25504 3927 25556 3936
rect 25504 3893 25513 3927
rect 25513 3893 25547 3927
rect 25547 3893 25556 3927
rect 25504 3884 25556 3893
rect 28540 3884 28592 3936
rect 29460 3884 29512 3936
rect 37740 4088 37792 4140
rect 37188 3952 37240 4004
rect 37280 3927 37332 3936
rect 37280 3893 37289 3927
rect 37289 3893 37323 3927
rect 37323 3893 37332 3927
rect 37280 3884 37332 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 7472 3680 7524 3732
rect 7840 3723 7892 3732
rect 7840 3689 7849 3723
rect 7849 3689 7883 3723
rect 7883 3689 7892 3723
rect 7840 3680 7892 3689
rect 8760 3680 8812 3732
rect 9588 3680 9640 3732
rect 10232 3680 10284 3732
rect 13452 3680 13504 3732
rect 14372 3723 14424 3732
rect 14372 3689 14381 3723
rect 14381 3689 14415 3723
rect 14415 3689 14424 3723
rect 14372 3680 14424 3689
rect 16580 3680 16632 3732
rect 17132 3680 17184 3732
rect 18420 3680 18472 3732
rect 18880 3680 18932 3732
rect 19340 3680 19392 3732
rect 22744 3723 22796 3732
rect 6184 3655 6236 3664
rect 6184 3621 6193 3655
rect 6193 3621 6227 3655
rect 6227 3621 6236 3655
rect 6184 3612 6236 3621
rect 12624 3612 12676 3664
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 8208 3476 8260 3528
rect 9588 3476 9640 3528
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 11704 3544 11756 3596
rect 12164 3587 12216 3596
rect 12164 3553 12173 3587
rect 12173 3553 12207 3587
rect 12207 3553 12216 3587
rect 12164 3544 12216 3553
rect 13268 3612 13320 3664
rect 15660 3612 15712 3664
rect 20720 3612 20772 3664
rect 21272 3612 21324 3664
rect 22744 3689 22753 3723
rect 22753 3689 22787 3723
rect 22787 3689 22796 3723
rect 22744 3680 22796 3689
rect 23020 3680 23072 3732
rect 26424 3680 26476 3732
rect 27068 3680 27120 3732
rect 29000 3723 29052 3732
rect 29000 3689 29009 3723
rect 29009 3689 29043 3723
rect 29043 3689 29052 3723
rect 29000 3680 29052 3689
rect 29092 3680 29144 3732
rect 30104 3723 30156 3732
rect 30104 3689 30113 3723
rect 30113 3689 30147 3723
rect 30147 3689 30156 3723
rect 30104 3680 30156 3689
rect 33600 3680 33652 3732
rect 28448 3612 28500 3664
rect 36544 3612 36596 3664
rect 38108 3612 38160 3664
rect 6828 3408 6880 3460
rect 6920 3408 6972 3460
rect 11152 3476 11204 3528
rect 11520 3519 11572 3528
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11520 3476 11572 3485
rect 12992 3544 13044 3596
rect 2872 3340 2924 3392
rect 4896 3340 4948 3392
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 10048 3340 10100 3392
rect 10876 3340 10928 3392
rect 11888 3408 11940 3460
rect 12532 3485 12541 3506
rect 12541 3485 12575 3506
rect 12575 3485 12584 3506
rect 12532 3454 12584 3485
rect 12900 3476 12952 3528
rect 14556 3544 14608 3596
rect 14832 3544 14884 3596
rect 16488 3587 16540 3596
rect 16488 3553 16497 3587
rect 16497 3553 16531 3587
rect 16531 3553 16540 3587
rect 16488 3544 16540 3553
rect 16856 3544 16908 3596
rect 19708 3587 19760 3596
rect 19708 3553 19717 3587
rect 19717 3553 19751 3587
rect 19751 3553 19760 3587
rect 19708 3544 19760 3553
rect 20168 3544 20220 3596
rect 21088 3544 21140 3596
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 16396 3519 16448 3528
rect 14280 3408 14332 3460
rect 15108 3451 15160 3460
rect 15108 3417 15117 3451
rect 15117 3417 15151 3451
rect 15151 3417 15160 3451
rect 15108 3408 15160 3417
rect 12532 3340 12584 3392
rect 13728 3340 13780 3392
rect 13820 3340 13872 3392
rect 15292 3340 15344 3392
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16396 3476 16448 3485
rect 16764 3476 16816 3528
rect 20536 3476 20588 3528
rect 21180 3476 21232 3528
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21364 3476 21416 3485
rect 23848 3476 23900 3528
rect 24584 3476 24636 3528
rect 26240 3544 26292 3596
rect 26424 3544 26476 3596
rect 26884 3544 26936 3596
rect 27160 3544 27212 3596
rect 24768 3476 24820 3528
rect 16672 3451 16724 3460
rect 16672 3417 16681 3451
rect 16681 3417 16715 3451
rect 16715 3417 16724 3451
rect 16672 3408 16724 3417
rect 23940 3408 23992 3460
rect 16304 3340 16356 3392
rect 20076 3340 20128 3392
rect 22836 3340 22888 3392
rect 23848 3340 23900 3392
rect 24952 3340 25004 3392
rect 25596 3476 25648 3528
rect 27804 3519 27856 3528
rect 27804 3485 27813 3519
rect 27813 3485 27847 3519
rect 27847 3485 27856 3519
rect 27804 3476 27856 3485
rect 33048 3544 33100 3596
rect 36360 3587 36412 3596
rect 36360 3553 36369 3587
rect 36369 3553 36403 3587
rect 36403 3553 36412 3587
rect 36360 3544 36412 3553
rect 33784 3476 33836 3528
rect 35348 3476 35400 3528
rect 37740 3544 37792 3596
rect 37004 3519 37056 3528
rect 37004 3485 37013 3519
rect 37013 3485 37047 3519
rect 37047 3485 37056 3519
rect 37004 3476 37056 3485
rect 37648 3519 37700 3528
rect 37648 3485 37657 3519
rect 37657 3485 37691 3519
rect 37691 3485 37700 3519
rect 37648 3476 37700 3485
rect 32220 3408 32272 3460
rect 35992 3408 36044 3460
rect 37556 3408 37608 3460
rect 28448 3340 28500 3392
rect 30196 3340 30248 3392
rect 31484 3383 31536 3392
rect 31484 3349 31493 3383
rect 31493 3349 31527 3383
rect 31527 3349 31536 3383
rect 31484 3340 31536 3349
rect 33416 3340 33468 3392
rect 33600 3340 33652 3392
rect 33784 3383 33836 3392
rect 33784 3349 33793 3383
rect 33793 3349 33827 3383
rect 33827 3349 33836 3383
rect 33784 3340 33836 3349
rect 34796 3340 34848 3392
rect 35808 3340 35860 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 5816 3179 5868 3188
rect 5816 3145 5825 3179
rect 5825 3145 5859 3179
rect 5859 3145 5868 3179
rect 5816 3136 5868 3145
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 9588 3179 9640 3188
rect 9588 3145 9597 3179
rect 9597 3145 9631 3179
rect 9631 3145 9640 3179
rect 9588 3136 9640 3145
rect 12532 3136 12584 3188
rect 13636 3136 13688 3188
rect 15108 3136 15160 3188
rect 15936 3179 15988 3188
rect 6920 3068 6972 3120
rect 9036 3068 9088 3120
rect 4620 3000 4672 3052
rect 5080 3000 5132 3052
rect 5264 3000 5316 3052
rect 5632 3043 5684 3052
rect 5632 3009 5641 3043
rect 5641 3009 5675 3043
rect 5675 3009 5684 3043
rect 5632 3000 5684 3009
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 7840 3000 7892 3052
rect 8116 3000 8168 3052
rect 8852 3000 8904 3052
rect 10048 3000 10100 3052
rect 10232 3043 10284 3052
rect 10232 3009 10241 3043
rect 10241 3009 10275 3043
rect 10275 3009 10284 3043
rect 10232 3000 10284 3009
rect 10692 3000 10744 3052
rect 9128 2975 9180 2984
rect 9128 2941 9137 2975
rect 9137 2941 9171 2975
rect 9171 2941 9180 2975
rect 9128 2932 9180 2941
rect 11888 3068 11940 3120
rect 15936 3145 15945 3179
rect 15945 3145 15979 3179
rect 15979 3145 15988 3179
rect 15936 3136 15988 3145
rect 17408 3179 17460 3188
rect 17408 3145 17417 3179
rect 17417 3145 17451 3179
rect 17451 3145 17460 3179
rect 17408 3136 17460 3145
rect 17592 3136 17644 3188
rect 19984 3179 20036 3188
rect 19984 3145 19993 3179
rect 19993 3145 20027 3179
rect 20027 3145 20036 3179
rect 19984 3136 20036 3145
rect 19340 3068 19392 3120
rect 11796 3000 11848 3052
rect 9956 2864 10008 2916
rect 10876 2932 10928 2984
rect 11888 2975 11940 2984
rect 11888 2941 11897 2975
rect 11897 2941 11931 2975
rect 11931 2941 11940 2975
rect 11888 2932 11940 2941
rect 12808 2932 12860 2984
rect 1768 2839 1820 2848
rect 1768 2805 1777 2839
rect 1777 2805 1811 2839
rect 1811 2805 1820 2839
rect 1768 2796 1820 2805
rect 2320 2839 2372 2848
rect 2320 2805 2329 2839
rect 2329 2805 2363 2839
rect 2363 2805 2372 2839
rect 2320 2796 2372 2805
rect 3424 2796 3476 2848
rect 5172 2839 5224 2848
rect 5172 2805 5181 2839
rect 5181 2805 5215 2839
rect 5215 2805 5224 2839
rect 5172 2796 5224 2805
rect 8392 2839 8444 2848
rect 8392 2805 8401 2839
rect 8401 2805 8435 2839
rect 8435 2805 8444 2839
rect 8392 2796 8444 2805
rect 13820 3000 13872 3052
rect 14004 3000 14056 3052
rect 13452 2932 13504 2984
rect 15108 2864 15160 2916
rect 13636 2839 13688 2848
rect 13636 2805 13645 2839
rect 13645 2805 13679 2839
rect 13679 2805 13688 2839
rect 13636 2796 13688 2805
rect 14740 2839 14792 2848
rect 14740 2805 14749 2839
rect 14749 2805 14783 2839
rect 14783 2805 14792 2839
rect 14740 2796 14792 2805
rect 15384 2932 15436 2984
rect 15752 3000 15804 3052
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 16948 3000 17000 3009
rect 17868 3000 17920 3052
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 16856 2975 16908 2984
rect 16856 2941 16865 2975
rect 16865 2941 16899 2975
rect 16899 2941 16908 2975
rect 16856 2932 16908 2941
rect 17500 2932 17552 2984
rect 18788 2932 18840 2984
rect 19340 2932 19392 2984
rect 20168 3068 20220 3120
rect 19616 3043 19668 3052
rect 19616 3009 19625 3043
rect 19625 3009 19659 3043
rect 19659 3009 19668 3043
rect 19616 3000 19668 3009
rect 20168 2932 20220 2984
rect 23020 3136 23072 3188
rect 23204 3179 23256 3188
rect 23204 3145 23213 3179
rect 23213 3145 23247 3179
rect 23247 3145 23256 3179
rect 23204 3136 23256 3145
rect 24032 3136 24084 3188
rect 25872 3179 25924 3188
rect 20996 3000 21048 3052
rect 21364 3000 21416 3052
rect 23480 3068 23532 3120
rect 24124 3068 24176 3120
rect 25872 3145 25881 3179
rect 25881 3145 25915 3179
rect 25915 3145 25924 3179
rect 25872 3136 25924 3145
rect 30840 3179 30892 3188
rect 30840 3145 30849 3179
rect 30849 3145 30883 3179
rect 30883 3145 30892 3179
rect 30840 3136 30892 3145
rect 33784 3136 33836 3188
rect 33968 3179 34020 3188
rect 33968 3145 33977 3179
rect 33977 3145 34011 3179
rect 34011 3145 34020 3179
rect 33968 3136 34020 3145
rect 35716 3136 35768 3188
rect 35992 3136 36044 3188
rect 37924 3136 37976 3188
rect 22100 3043 22152 3052
rect 22100 3009 22134 3043
rect 22134 3009 22152 3043
rect 22100 3000 22152 3009
rect 16120 2796 16172 2848
rect 18604 2796 18656 2848
rect 20168 2796 20220 2848
rect 20536 2796 20588 2848
rect 22192 2796 22244 2848
rect 24584 3000 24636 3052
rect 27436 3068 27488 3120
rect 28080 3111 28132 3120
rect 28080 3077 28098 3111
rect 28098 3077 28132 3111
rect 28080 3068 28132 3077
rect 29644 3068 29696 3120
rect 30196 3068 30248 3120
rect 28356 3043 28408 3052
rect 28356 3009 28365 3043
rect 28365 3009 28399 3043
rect 28399 3009 28408 3043
rect 28356 3000 28408 3009
rect 30104 3000 30156 3052
rect 30564 3000 30616 3052
rect 31024 3000 31076 3052
rect 32772 3068 32824 3120
rect 37280 3068 37332 3120
rect 37648 3068 37700 3120
rect 38016 3111 38068 3120
rect 38016 3077 38025 3111
rect 38025 3077 38059 3111
rect 38059 3077 38068 3111
rect 38016 3068 38068 3077
rect 31760 3000 31812 3052
rect 34152 3043 34204 3052
rect 34152 3009 34161 3043
rect 34161 3009 34195 3043
rect 34195 3009 34204 3043
rect 34152 3000 34204 3009
rect 36360 3000 36412 3052
rect 31484 2932 31536 2984
rect 32128 2975 32180 2984
rect 32128 2941 32137 2975
rect 32137 2941 32171 2975
rect 32171 2941 32180 2975
rect 32128 2932 32180 2941
rect 26884 2864 26936 2916
rect 29460 2796 29512 2848
rect 31300 2864 31352 2916
rect 30472 2796 30524 2848
rect 33508 2839 33560 2848
rect 33508 2805 33517 2839
rect 33517 2805 33551 2839
rect 33551 2805 33560 2839
rect 33508 2796 33560 2805
rect 34336 2796 34388 2848
rect 37556 2796 37608 2848
rect 38292 2796 38344 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 8668 2592 8720 2644
rect 7472 2456 7524 2508
rect 1768 2388 1820 2440
rect 2320 2388 2372 2440
rect 2872 2388 2924 2440
rect 5540 2388 5592 2440
rect 7288 2388 7340 2440
rect 8208 2431 8260 2440
rect 5724 2320 5776 2372
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 9680 2592 9732 2644
rect 9956 2592 10008 2644
rect 11888 2592 11940 2644
rect 12348 2592 12400 2644
rect 14556 2592 14608 2644
rect 14832 2635 14884 2644
rect 14832 2601 14841 2635
rect 14841 2601 14875 2635
rect 14875 2601 14884 2635
rect 14832 2592 14884 2601
rect 16856 2592 16908 2644
rect 18328 2592 18380 2644
rect 19432 2592 19484 2644
rect 20444 2635 20496 2644
rect 20444 2601 20453 2635
rect 20453 2601 20487 2635
rect 20487 2601 20496 2635
rect 20444 2592 20496 2601
rect 11796 2524 11848 2576
rect 12256 2524 12308 2576
rect 26516 2592 26568 2644
rect 26608 2592 26660 2644
rect 30656 2592 30708 2644
rect 31668 2592 31720 2644
rect 11060 2456 11112 2508
rect 8484 2388 8536 2440
rect 9036 2431 9088 2440
rect 9036 2397 9045 2431
rect 9045 2397 9079 2431
rect 9079 2397 9088 2431
rect 9036 2388 9088 2397
rect 9496 2388 9548 2440
rect 10508 2431 10560 2440
rect 8300 2320 8352 2372
rect 10508 2397 10517 2431
rect 10517 2397 10551 2431
rect 10551 2397 10560 2431
rect 10508 2388 10560 2397
rect 11152 2320 11204 2372
rect 1860 2295 1912 2304
rect 1860 2261 1869 2295
rect 1869 2261 1903 2295
rect 1903 2261 1912 2295
rect 1860 2252 1912 2261
rect 5172 2295 5224 2304
rect 5172 2261 5181 2295
rect 5181 2261 5215 2295
rect 5215 2261 5224 2295
rect 5172 2252 5224 2261
rect 5816 2295 5868 2304
rect 5816 2261 5825 2295
rect 5825 2261 5859 2295
rect 5859 2261 5868 2295
rect 5816 2252 5868 2261
rect 12440 2388 12492 2440
rect 12624 2388 12676 2440
rect 13452 2456 13504 2508
rect 15200 2456 15252 2508
rect 17224 2456 17276 2508
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 12348 2252 12400 2304
rect 14464 2320 14516 2372
rect 15016 2320 15068 2372
rect 16672 2388 16724 2440
rect 16948 2431 17000 2440
rect 16948 2397 16957 2431
rect 16957 2397 16991 2431
rect 16991 2397 17000 2431
rect 16948 2388 17000 2397
rect 19156 2456 19208 2508
rect 19340 2499 19392 2508
rect 19340 2465 19349 2499
rect 19349 2465 19383 2499
rect 19383 2465 19392 2499
rect 19340 2456 19392 2465
rect 20168 2456 20220 2508
rect 24400 2524 24452 2576
rect 24124 2456 24176 2508
rect 25504 2456 25556 2508
rect 29000 2524 29052 2576
rect 32496 2524 32548 2576
rect 33600 2592 33652 2644
rect 36452 2592 36504 2644
rect 13544 2295 13596 2304
rect 13544 2261 13553 2295
rect 13553 2261 13587 2295
rect 13587 2261 13596 2295
rect 13544 2252 13596 2261
rect 14188 2295 14240 2304
rect 14188 2261 14197 2295
rect 14197 2261 14231 2295
rect 14231 2261 14240 2295
rect 14188 2252 14240 2261
rect 17960 2388 18012 2440
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 18696 2388 18748 2440
rect 20720 2388 20772 2440
rect 22468 2388 22520 2440
rect 25044 2388 25096 2440
rect 18880 2320 18932 2372
rect 19616 2363 19668 2372
rect 19616 2329 19625 2363
rect 19625 2329 19659 2363
rect 19659 2329 19668 2363
rect 19616 2320 19668 2329
rect 20076 2320 20128 2372
rect 26332 2388 26384 2440
rect 28724 2431 28776 2440
rect 17960 2252 18012 2304
rect 18512 2252 18564 2304
rect 19432 2252 19484 2304
rect 21088 2295 21140 2304
rect 21088 2261 21097 2295
rect 21097 2261 21131 2295
rect 21131 2261 21140 2295
rect 21088 2252 21140 2261
rect 23296 2252 23348 2304
rect 24492 2295 24544 2304
rect 24492 2261 24501 2295
rect 24501 2261 24535 2295
rect 24535 2261 24544 2295
rect 24492 2252 24544 2261
rect 26056 2252 26108 2304
rect 28724 2397 28733 2431
rect 28733 2397 28767 2431
rect 28767 2397 28776 2431
rect 28724 2388 28776 2397
rect 28080 2320 28132 2372
rect 29368 2388 29420 2440
rect 29000 2320 29052 2372
rect 29828 2320 29880 2372
rect 31300 2388 31352 2440
rect 32128 2456 32180 2508
rect 37556 2499 37608 2508
rect 37556 2465 37565 2499
rect 37565 2465 37599 2499
rect 37599 2465 37608 2499
rect 37556 2456 37608 2465
rect 34244 2388 34296 2440
rect 34796 2388 34848 2440
rect 36636 2388 36688 2440
rect 37096 2388 37148 2440
rect 37832 2388 37884 2440
rect 29092 2252 29144 2304
rect 29552 2295 29604 2304
rect 29552 2261 29561 2295
rect 29561 2261 29595 2295
rect 29595 2261 29604 2295
rect 29552 2252 29604 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 1860 2048 1912 2100
rect 5816 2048 5868 2100
rect 9864 2048 9916 2100
rect 10968 2048 11020 2100
rect 13452 2048 13504 2100
rect 13544 2048 13596 2100
rect 16580 2048 16632 2100
rect 21640 2048 21692 2100
rect 24492 2048 24544 2100
rect 26516 2048 26568 2100
rect 29644 2048 29696 2100
rect 8760 1980 8812 2032
rect 14188 1980 14240 2032
rect 18420 1980 18472 2032
rect 5724 1912 5776 1964
rect 8576 1912 8628 1964
rect 17868 1912 17920 1964
rect 29552 1912 29604 1964
rect 5172 1844 5224 1896
rect 12440 1844 12492 1896
rect 13360 1844 13412 1896
rect 13728 1844 13780 1896
rect 20076 1844 20128 1896
rect 11612 1776 11664 1828
rect 16948 1776 17000 1828
rect 5540 1708 5592 1760
rect 6184 1708 6236 1760
rect 8208 1708 8260 1760
rect 9496 1708 9548 1760
rect 12624 1708 12676 1760
rect 14464 1708 14516 1760
rect 16856 1368 16908 1420
rect 17776 1368 17828 1420
<< metal2 >>
rect 1766 39200 1822 40000
rect 2318 39200 2374 40000
rect 2870 39200 2926 40000
rect 3422 39200 3478 40000
rect 3974 39200 4030 40000
rect 4526 39200 4582 40000
rect 5078 39200 5134 40000
rect 5630 39200 5686 40000
rect 6182 39200 6238 40000
rect 6734 39200 6790 40000
rect 7286 39200 7342 40000
rect 7838 39200 7894 40000
rect 8390 39200 8446 40000
rect 8942 39200 8998 40000
rect 9494 39200 9550 40000
rect 10046 39200 10102 40000
rect 10598 39200 10654 40000
rect 11150 39200 11206 40000
rect 11702 39200 11758 40000
rect 12254 39200 12310 40000
rect 12806 39200 12862 40000
rect 13358 39200 13414 40000
rect 13910 39200 13966 40000
rect 14462 39200 14518 40000
rect 15014 39200 15070 40000
rect 15566 39200 15622 40000
rect 16118 39200 16174 40000
rect 16670 39200 16726 40000
rect 17222 39200 17278 40000
rect 17774 39200 17830 40000
rect 17972 39222 18276 39250
rect 1780 37262 1808 39200
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 1780 36922 1808 37198
rect 2332 37126 2360 39200
rect 2504 37256 2556 37262
rect 2504 37198 2556 37204
rect 2320 37120 2372 37126
rect 2320 37062 2372 37068
rect 1768 36916 1820 36922
rect 1768 36858 1820 36864
rect 2516 36242 2544 37198
rect 2884 37126 2912 39200
rect 3240 37256 3292 37262
rect 3240 37198 3292 37204
rect 2872 37120 2924 37126
rect 2872 37062 2924 37068
rect 3252 36922 3280 37198
rect 3240 36916 3292 36922
rect 3240 36858 3292 36864
rect 3436 36854 3464 39200
rect 3988 37108 4016 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4160 37120 4212 37126
rect 3988 37080 4160 37108
rect 4160 37062 4212 37068
rect 4632 36922 4660 37726
rect 4712 37256 4764 37262
rect 4712 37198 4764 37204
rect 4620 36916 4672 36922
rect 4620 36858 4672 36864
rect 3424 36848 3476 36854
rect 3424 36790 3476 36796
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 2504 36236 2556 36242
rect 2504 36178 2556 36184
rect 4724 36038 4752 37198
rect 5092 37126 5120 39200
rect 5644 37126 5672 39200
rect 5816 37256 5868 37262
rect 5816 37198 5868 37204
rect 5080 37120 5132 37126
rect 5080 37062 5132 37068
rect 5632 37120 5684 37126
rect 5632 37062 5684 37068
rect 5080 36780 5132 36786
rect 5080 36722 5132 36728
rect 5092 36038 5120 36722
rect 5828 36582 5856 37198
rect 6196 36922 6224 39200
rect 6748 37126 6776 39200
rect 7012 37188 7064 37194
rect 7012 37130 7064 37136
rect 6736 37120 6788 37126
rect 6736 37062 6788 37068
rect 6184 36916 6236 36922
rect 6184 36858 6236 36864
rect 6644 36780 6696 36786
rect 6644 36722 6696 36728
rect 5816 36576 5868 36582
rect 5816 36518 5868 36524
rect 4712 36032 4764 36038
rect 4712 35974 4764 35980
rect 5080 36032 5132 36038
rect 5080 35974 5132 35980
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4724 31210 4752 35974
rect 5092 32502 5120 35974
rect 5080 32496 5132 32502
rect 5080 32438 5132 32444
rect 4712 31204 4764 31210
rect 4712 31146 4764 31152
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5828 28558 5856 36518
rect 6656 36310 6684 36722
rect 6828 36644 6880 36650
rect 6828 36586 6880 36592
rect 6644 36304 6696 36310
rect 6644 36246 6696 36252
rect 6840 35086 6868 36586
rect 7024 36106 7052 37130
rect 7300 37126 7328 39200
rect 7380 37256 7432 37262
rect 7380 37198 7432 37204
rect 7288 37120 7340 37126
rect 7288 37062 7340 37068
rect 7392 36582 7420 37198
rect 7852 36922 7880 39200
rect 8300 37188 8352 37194
rect 8300 37130 8352 37136
rect 7840 36916 7892 36922
rect 7840 36858 7892 36864
rect 8208 36780 8260 36786
rect 8208 36722 8260 36728
rect 7380 36576 7432 36582
rect 7380 36518 7432 36524
rect 7012 36100 7064 36106
rect 7012 36042 7064 36048
rect 6828 35080 6880 35086
rect 6828 35022 6880 35028
rect 5816 28552 5868 28558
rect 5816 28494 5868 28500
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 7392 26382 7420 36518
rect 7564 36100 7616 36106
rect 7564 36042 7616 36048
rect 7576 27334 7604 36042
rect 8220 36038 8248 36722
rect 8312 36174 8340 37130
rect 8404 37126 8432 39200
rect 8576 37256 8628 37262
rect 8576 37198 8628 37204
rect 8392 37120 8444 37126
rect 8392 37062 8444 37068
rect 8300 36168 8352 36174
rect 8300 36110 8352 36116
rect 8208 36032 8260 36038
rect 8208 35974 8260 35980
rect 8588 35494 8616 37198
rect 8956 36922 8984 39200
rect 9508 37126 9536 39200
rect 9956 37392 10008 37398
rect 9956 37334 10008 37340
rect 9496 37120 9548 37126
rect 9496 37062 9548 37068
rect 8944 36916 8996 36922
rect 8944 36858 8996 36864
rect 9680 36848 9732 36854
rect 9680 36790 9732 36796
rect 9312 36780 9364 36786
rect 9312 36722 9364 36728
rect 9324 36242 9352 36722
rect 8760 36236 8812 36242
rect 8760 36178 8812 36184
rect 9312 36236 9364 36242
rect 9312 36178 9364 36184
rect 8576 35488 8628 35494
rect 8576 35430 8628 35436
rect 8588 29102 8616 35430
rect 8772 33658 8800 36178
rect 8944 36168 8996 36174
rect 8944 36110 8996 36116
rect 8760 33652 8812 33658
rect 8760 33594 8812 33600
rect 8852 33516 8904 33522
rect 8852 33458 8904 33464
rect 8576 29096 8628 29102
rect 8576 29038 8628 29044
rect 7564 27328 7616 27334
rect 7564 27270 7616 27276
rect 8576 26988 8628 26994
rect 8576 26930 8628 26936
rect 7380 26376 7432 26382
rect 7380 26318 7432 26324
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 8588 25498 8616 26930
rect 8760 26784 8812 26790
rect 8760 26726 8812 26732
rect 8772 25906 8800 26726
rect 8760 25900 8812 25906
rect 8760 25842 8812 25848
rect 8576 25492 8628 25498
rect 8576 25434 8628 25440
rect 8864 25265 8892 33458
rect 8956 25362 8984 36110
rect 9692 34950 9720 36790
rect 9680 34944 9732 34950
rect 9680 34886 9732 34892
rect 9404 34740 9456 34746
rect 9404 34682 9456 34688
rect 9416 33998 9444 34682
rect 9220 33992 9272 33998
rect 9220 33934 9272 33940
rect 9404 33992 9456 33998
rect 9404 33934 9456 33940
rect 9232 33454 9260 33934
rect 9692 33522 9720 34886
rect 9968 34678 9996 37334
rect 10060 37126 10088 39200
rect 10324 37256 10376 37262
rect 10244 37216 10324 37244
rect 10048 37120 10100 37126
rect 10048 37062 10100 37068
rect 10244 36582 10272 37216
rect 10324 37198 10376 37204
rect 10416 37188 10468 37194
rect 10416 37130 10468 37136
rect 10232 36576 10284 36582
rect 10232 36518 10284 36524
rect 10048 36304 10100 36310
rect 10048 36246 10100 36252
rect 9956 34672 10008 34678
rect 9956 34614 10008 34620
rect 9680 33516 9732 33522
rect 9680 33458 9732 33464
rect 9220 33448 9272 33454
rect 9220 33390 9272 33396
rect 9692 33114 9720 33458
rect 9680 33108 9732 33114
rect 9680 33050 9732 33056
rect 10060 31754 10088 36246
rect 10244 36145 10272 36518
rect 10428 36174 10456 37130
rect 10612 36922 10640 39200
rect 11060 37188 11112 37194
rect 11060 37130 11112 37136
rect 10600 36916 10652 36922
rect 10600 36858 10652 36864
rect 10968 36780 11020 36786
rect 10968 36722 11020 36728
rect 10416 36168 10468 36174
rect 10230 36136 10286 36145
rect 10416 36110 10468 36116
rect 10980 36106 11008 36722
rect 10230 36071 10286 36080
rect 10968 36100 11020 36106
rect 10968 36042 11020 36048
rect 11072 35494 11100 37130
rect 11164 37126 11192 39200
rect 11716 37126 11744 39200
rect 12072 37256 12124 37262
rect 12072 37198 12124 37204
rect 11152 37120 11204 37126
rect 11152 37062 11204 37068
rect 11704 37120 11756 37126
rect 11704 37062 11756 37068
rect 12084 36038 12112 37198
rect 12268 36904 12296 39200
rect 12532 37256 12584 37262
rect 12532 37198 12584 37204
rect 12440 36916 12492 36922
rect 12268 36876 12440 36904
rect 12440 36858 12492 36864
rect 12544 36582 12572 37198
rect 12820 37126 12848 39200
rect 13372 37126 13400 39200
rect 13452 37664 13504 37670
rect 13452 37606 13504 37612
rect 12808 37120 12860 37126
rect 12808 37062 12860 37068
rect 13360 37120 13412 37126
rect 13360 37062 13412 37068
rect 12624 36780 12676 36786
rect 12624 36722 12676 36728
rect 12532 36576 12584 36582
rect 12532 36518 12584 36524
rect 11428 36032 11480 36038
rect 11428 35974 11480 35980
rect 12072 36032 12124 36038
rect 12072 35974 12124 35980
rect 11060 35488 11112 35494
rect 11060 35430 11112 35436
rect 10876 35284 10928 35290
rect 10876 35226 10928 35232
rect 10140 35012 10192 35018
rect 10140 34954 10192 34960
rect 10152 34542 10180 34954
rect 10888 34746 10916 35226
rect 10876 34740 10928 34746
rect 10876 34682 10928 34688
rect 10232 34604 10284 34610
rect 10232 34546 10284 34552
rect 10324 34604 10376 34610
rect 10324 34546 10376 34552
rect 10140 34536 10192 34542
rect 10140 34478 10192 34484
rect 10244 33998 10272 34546
rect 10336 34202 10364 34546
rect 10324 34196 10376 34202
rect 10324 34138 10376 34144
rect 10232 33992 10284 33998
rect 10232 33934 10284 33940
rect 10244 33658 10272 33934
rect 10232 33652 10284 33658
rect 10232 33594 10284 33600
rect 10060 31726 10180 31754
rect 10152 29578 10180 31726
rect 10140 29572 10192 29578
rect 10140 29514 10192 29520
rect 10152 29306 10180 29514
rect 10140 29300 10192 29306
rect 10140 29242 10192 29248
rect 9588 28960 9640 28966
rect 9588 28902 9640 28908
rect 9600 28626 9628 28902
rect 9588 28620 9640 28626
rect 9588 28562 9640 28568
rect 9128 28552 9180 28558
rect 9128 28494 9180 28500
rect 9036 28416 9088 28422
rect 9036 28358 9088 28364
rect 9048 28082 9076 28358
rect 9036 28076 9088 28082
rect 9036 28018 9088 28024
rect 9140 27962 9168 28494
rect 9048 27934 9168 27962
rect 8944 25356 8996 25362
rect 8944 25298 8996 25304
rect 8850 25256 8906 25265
rect 8850 25191 8906 25200
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 9048 9654 9076 27934
rect 9494 27432 9550 27441
rect 9494 27367 9550 27376
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 9140 26586 9168 26930
rect 9128 26580 9180 26586
rect 9128 26522 9180 26528
rect 9508 26042 9536 27367
rect 9600 26450 9628 28562
rect 10152 28506 10180 29242
rect 10508 29028 10560 29034
rect 10508 28970 10560 28976
rect 10520 28558 10548 28970
rect 10876 28960 10928 28966
rect 10876 28902 10928 28908
rect 10888 28558 10916 28902
rect 10060 28478 10180 28506
rect 10508 28552 10560 28558
rect 10508 28494 10560 28500
rect 10876 28552 10928 28558
rect 10876 28494 10928 28500
rect 10060 28422 10088 28478
rect 10048 28416 10100 28422
rect 10048 28358 10100 28364
rect 10232 28416 10284 28422
rect 10232 28358 10284 28364
rect 9956 28212 10008 28218
rect 9956 28154 10008 28160
rect 9968 28121 9996 28154
rect 9954 28112 10010 28121
rect 10244 28082 10272 28358
rect 9954 28047 10010 28056
rect 10232 28076 10284 28082
rect 10232 28018 10284 28024
rect 10508 27396 10560 27402
rect 10508 27338 10560 27344
rect 10230 26888 10286 26897
rect 10230 26823 10232 26832
rect 10284 26823 10286 26832
rect 10232 26794 10284 26800
rect 9588 26444 9640 26450
rect 9588 26386 9640 26392
rect 9864 26308 9916 26314
rect 9864 26250 9916 26256
rect 9496 26036 9548 26042
rect 9496 25978 9548 25984
rect 9876 25702 9904 26250
rect 9864 25696 9916 25702
rect 9864 25638 9916 25644
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 9600 24954 9628 25298
rect 9588 24948 9640 24954
rect 9588 24890 9640 24896
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9036 9648 9088 9654
rect 9036 9590 9088 9596
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4080 3534 4108 3878
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 1780 2446 1808 2790
rect 2332 2446 2360 2790
rect 2884 2446 2912 3334
rect 3424 2848 3476 2854
rect 3424 2790 3476 2796
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 1780 800 1808 2382
rect 1860 2304 1912 2310
rect 1860 2246 1912 2252
rect 1872 2106 1900 2246
rect 1860 2100 1912 2106
rect 1860 2042 1912 2048
rect 2332 800 2360 2382
rect 2884 800 2912 2382
rect 3436 800 3464 2790
rect 4080 2774 4108 3470
rect 4632 3058 4660 3878
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 3988 2746 4108 2774
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 3988 800 4016 2746
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 1442 4660 2994
rect 4908 2774 4936 3334
rect 5276 3058 5304 4422
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 4908 2746 5028 2774
rect 5000 2417 5028 2746
rect 4986 2408 5042 2417
rect 4986 2343 5042 2352
rect 4540 1414 4660 1442
rect 4540 800 4568 1414
rect 5092 800 5120 2994
rect 5170 2952 5226 2961
rect 5170 2887 5226 2896
rect 5184 2854 5212 2887
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5552 2446 5580 3878
rect 5644 3058 5672 4422
rect 5828 3194 5856 9522
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 6184 3664 6236 3670
rect 6182 3632 6184 3641
rect 6236 3632 6238 3641
rect 6182 3567 6238 3576
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6840 3058 6868 3402
rect 6932 3126 6960 3402
rect 7024 3194 7052 7414
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7208 3777 7236 3878
rect 7194 3768 7250 3777
rect 7194 3703 7250 3712
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5184 1902 5212 2246
rect 5172 1896 5224 1902
rect 5172 1838 5224 1844
rect 5552 1766 5580 2382
rect 5540 1760 5592 1766
rect 5540 1702 5592 1708
rect 5644 800 5672 2994
rect 6840 2774 6868 2994
rect 6748 2746 6868 2774
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5736 1970 5764 2314
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5828 2106 5856 2246
rect 5816 2100 5868 2106
rect 5816 2042 5868 2048
rect 5724 1964 5776 1970
rect 5724 1906 5776 1912
rect 6184 1760 6236 1766
rect 6184 1702 6236 1708
rect 6196 800 6224 1702
rect 6748 800 6776 2746
rect 7300 2446 7328 3946
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7484 2514 7512 3674
rect 7576 3058 7604 4966
rect 7852 3738 7880 5034
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 8128 3058 8156 4490
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7300 800 7328 2382
rect 7852 800 7880 2994
rect 8220 2446 8248 3470
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8220 1766 8248 2382
rect 8312 2378 8340 5510
rect 8404 2854 8432 6326
rect 8484 5636 8536 5642
rect 8484 5578 8536 5584
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8496 2446 8524 5578
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 8208 1760 8260 1766
rect 8312 1748 8340 2314
rect 8588 1970 8616 4218
rect 8680 2650 8708 8502
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8772 2038 8800 3674
rect 9048 3126 9076 4014
rect 9140 3641 9168 24006
rect 9876 16574 9904 25638
rect 10232 25424 10284 25430
rect 10230 25392 10232 25401
rect 10284 25392 10286 25401
rect 10230 25327 10286 25336
rect 10416 25152 10468 25158
rect 10416 25094 10468 25100
rect 10428 16574 10456 25094
rect 9692 16546 9904 16574
rect 10336 16546 10456 16574
rect 9692 6458 9720 16546
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10244 9042 10272 9590
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10244 8945 10272 8978
rect 10230 8936 10286 8945
rect 9864 8900 9916 8906
rect 10230 8871 10286 8880
rect 9864 8842 9916 8848
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9692 5778 9720 6394
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9692 5681 9720 5714
rect 9678 5672 9734 5681
rect 9678 5607 9734 5616
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9404 4752 9456 4758
rect 9404 4694 9456 4700
rect 9416 4282 9444 4694
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9404 3936 9456 3942
rect 9402 3904 9404 3913
rect 9456 3904 9458 3913
rect 9402 3839 9458 3848
rect 9126 3632 9182 3641
rect 9126 3567 9182 3576
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8864 2774 8892 2994
rect 8864 2746 8984 2774
rect 8760 2032 8812 2038
rect 8760 1974 8812 1980
rect 8576 1964 8628 1970
rect 8576 1906 8628 1912
rect 8312 1720 8432 1748
rect 8208 1702 8260 1708
rect 8404 800 8432 1720
rect 8956 800 8984 2746
rect 9048 2446 9076 3062
rect 9140 2990 9168 3567
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9324 2009 9352 3334
rect 9508 2446 9536 4558
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9600 3738 9628 3878
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9600 3194 9628 3470
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9692 2650 9720 5170
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9876 2106 9904 8842
rect 10336 8090 10364 16546
rect 10416 9104 10468 9110
rect 10416 9046 10468 9052
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10336 7546 10364 8026
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9968 5914 9996 7346
rect 10428 7342 10456 9046
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10428 6390 10456 7278
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 10428 5710 10456 6326
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10060 4078 10088 5102
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 10060 3398 10088 4014
rect 10152 3534 10180 4626
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10244 3738 10272 4082
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10336 3618 10364 5238
rect 10428 5166 10456 5646
rect 10520 5370 10548 27338
rect 10888 26234 10916 28494
rect 11072 28098 11100 35430
rect 11072 28070 11192 28098
rect 11060 28008 11112 28014
rect 11060 27950 11112 27956
rect 11072 27674 11100 27950
rect 11060 27668 11112 27674
rect 11060 27610 11112 27616
rect 11072 27554 11100 27610
rect 10980 27526 11100 27554
rect 10980 26926 11008 27526
rect 11164 27470 11192 28070
rect 11060 27464 11112 27470
rect 11060 27406 11112 27412
rect 11152 27464 11204 27470
rect 11152 27406 11204 27412
rect 10968 26920 11020 26926
rect 10968 26862 11020 26868
rect 10980 26450 11008 26862
rect 10968 26444 11020 26450
rect 10968 26386 11020 26392
rect 10888 26206 11008 26234
rect 10784 25696 10836 25702
rect 10784 25638 10836 25644
rect 10796 24954 10824 25638
rect 10784 24948 10836 24954
rect 10784 24890 10836 24896
rect 10980 22166 11008 26206
rect 11072 25498 11100 27406
rect 11244 26988 11296 26994
rect 11244 26930 11296 26936
rect 11256 26586 11284 26930
rect 11244 26580 11296 26586
rect 11244 26522 11296 26528
rect 11060 25492 11112 25498
rect 11060 25434 11112 25440
rect 11440 24886 11468 35974
rect 11888 35624 11940 35630
rect 11888 35566 11940 35572
rect 11704 34944 11756 34950
rect 11704 34886 11756 34892
rect 11612 28552 11664 28558
rect 11612 28494 11664 28500
rect 11624 27674 11652 28494
rect 11716 27962 11744 34886
rect 11900 34678 11928 35566
rect 11888 34672 11940 34678
rect 12084 34649 12112 35974
rect 12438 35320 12494 35329
rect 12438 35255 12494 35264
rect 12452 35018 12480 35255
rect 12440 35012 12492 35018
rect 12440 34954 12492 34960
rect 12164 34944 12216 34950
rect 12164 34886 12216 34892
rect 11888 34614 11940 34620
rect 12070 34640 12126 34649
rect 11900 33998 11928 34614
rect 12176 34610 12204 34886
rect 12070 34575 12126 34584
rect 12164 34604 12216 34610
rect 11888 33992 11940 33998
rect 11888 33934 11940 33940
rect 11796 30728 11848 30734
rect 11796 30670 11848 30676
rect 11980 30728 12032 30734
rect 11980 30670 12032 30676
rect 11808 30190 11836 30670
rect 11796 30184 11848 30190
rect 11796 30126 11848 30132
rect 11808 28506 11836 30126
rect 11992 29850 12020 30670
rect 11980 29844 12032 29850
rect 11980 29786 12032 29792
rect 12084 28694 12112 34575
rect 12164 34546 12216 34552
rect 12348 34604 12400 34610
rect 12348 34546 12400 34552
rect 12254 34232 12310 34241
rect 12254 34167 12310 34176
rect 12268 34134 12296 34167
rect 12256 34128 12308 34134
rect 12256 34070 12308 34076
rect 12360 33114 12388 34546
rect 12348 33108 12400 33114
rect 12348 33050 12400 33056
rect 12256 32428 12308 32434
rect 12256 32370 12308 32376
rect 12268 30938 12296 32370
rect 12544 31754 12572 36518
rect 12636 36038 12664 36722
rect 12716 36236 12768 36242
rect 12716 36178 12768 36184
rect 12624 36032 12676 36038
rect 12624 35974 12676 35980
rect 12728 33402 12756 36178
rect 13176 36168 13228 36174
rect 13176 36110 13228 36116
rect 12900 35148 12952 35154
rect 12900 35090 12952 35096
rect 12912 34610 12940 35090
rect 12900 34604 12952 34610
rect 12900 34546 12952 34552
rect 12808 34536 12860 34542
rect 12808 34478 12860 34484
rect 12820 33522 12848 34478
rect 12912 33930 12940 34546
rect 13084 34468 13136 34474
rect 13084 34410 13136 34416
rect 12992 34400 13044 34406
rect 12992 34342 13044 34348
rect 13004 34066 13032 34342
rect 12992 34060 13044 34066
rect 12992 34002 13044 34008
rect 12900 33924 12952 33930
rect 12900 33866 12952 33872
rect 13096 33658 13124 34410
rect 13188 33658 13216 36110
rect 13268 36032 13320 36038
rect 13268 35974 13320 35980
rect 13084 33652 13136 33658
rect 13084 33594 13136 33600
rect 13176 33652 13228 33658
rect 13176 33594 13228 33600
rect 12808 33516 12860 33522
rect 12808 33458 12860 33464
rect 13176 33516 13228 33522
rect 13176 33458 13228 33464
rect 12728 33374 12848 33402
rect 12716 33312 12768 33318
rect 12716 33254 12768 33260
rect 12728 32910 12756 33254
rect 12716 32904 12768 32910
rect 12716 32846 12768 32852
rect 12452 31726 12572 31754
rect 12256 30932 12308 30938
rect 12256 30874 12308 30880
rect 12256 30252 12308 30258
rect 12256 30194 12308 30200
rect 12164 29164 12216 29170
rect 12164 29106 12216 29112
rect 12072 28688 12124 28694
rect 12072 28630 12124 28636
rect 11808 28478 11928 28506
rect 11796 28416 11848 28422
rect 11796 28358 11848 28364
rect 11808 28150 11836 28358
rect 11796 28144 11848 28150
rect 11796 28086 11848 28092
rect 11900 28082 11928 28478
rect 12176 28218 12204 29106
rect 12164 28212 12216 28218
rect 12164 28154 12216 28160
rect 11888 28076 11940 28082
rect 11888 28018 11940 28024
rect 12072 28076 12124 28082
rect 12072 28018 12124 28024
rect 11716 27934 11836 27962
rect 11704 27872 11756 27878
rect 11704 27814 11756 27820
rect 11612 27668 11664 27674
rect 11612 27610 11664 27616
rect 11716 26382 11744 27814
rect 11520 26376 11572 26382
rect 11520 26318 11572 26324
rect 11704 26376 11756 26382
rect 11704 26318 11756 26324
rect 11428 24880 11480 24886
rect 11428 24822 11480 24828
rect 11532 24682 11560 26318
rect 11520 24676 11572 24682
rect 11520 24618 11572 24624
rect 11808 23526 11836 27934
rect 12084 27674 12112 28018
rect 12072 27668 12124 27674
rect 12072 27610 12124 27616
rect 12268 27130 12296 30194
rect 12346 29064 12402 29073
rect 12346 28999 12348 29008
rect 12400 28999 12402 29008
rect 12348 28970 12400 28976
rect 12346 28520 12402 28529
rect 12346 28455 12348 28464
rect 12400 28455 12402 28464
rect 12348 28426 12400 28432
rect 12256 27124 12308 27130
rect 12256 27066 12308 27072
rect 11888 26512 11940 26518
rect 11888 26454 11940 26460
rect 11900 26353 11928 26454
rect 12256 26376 12308 26382
rect 11886 26344 11942 26353
rect 12256 26318 12308 26324
rect 11886 26279 11942 26288
rect 12164 25696 12216 25702
rect 12164 25638 12216 25644
rect 12176 25430 12204 25638
rect 12164 25424 12216 25430
rect 12164 25366 12216 25372
rect 12176 24750 12204 25366
rect 12268 25362 12296 26318
rect 12348 25696 12400 25702
rect 12348 25638 12400 25644
rect 12256 25356 12308 25362
rect 12256 25298 12308 25304
rect 12360 25158 12388 25638
rect 12452 25362 12480 31726
rect 12624 30728 12676 30734
rect 12624 30670 12676 30676
rect 12636 30326 12664 30670
rect 12624 30320 12676 30326
rect 12624 30262 12676 30268
rect 12624 30048 12676 30054
rect 12624 29990 12676 29996
rect 12636 29646 12664 29990
rect 12624 29640 12676 29646
rect 12624 29582 12676 29588
rect 12532 29096 12584 29102
rect 12532 29038 12584 29044
rect 12544 27130 12572 29038
rect 12532 27124 12584 27130
rect 12532 27066 12584 27072
rect 12440 25356 12492 25362
rect 12440 25298 12492 25304
rect 12348 25152 12400 25158
rect 12348 25094 12400 25100
rect 11980 24744 12032 24750
rect 11980 24686 12032 24692
rect 12164 24744 12216 24750
rect 12164 24686 12216 24692
rect 11992 24070 12020 24686
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 11796 23520 11848 23526
rect 11796 23462 11848 23468
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 11980 22160 12032 22166
rect 11980 22102 12032 22108
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 10874 10160 10930 10169
rect 10874 10095 10930 10104
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 8498 10732 8774
rect 10888 8634 10916 10095
rect 11532 9722 11560 10610
rect 11702 10568 11758 10577
rect 11702 10503 11704 10512
rect 11756 10503 11758 10512
rect 11704 10474 11756 10480
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11992 9654 12020 22102
rect 12360 12434 12388 25094
rect 12636 12434 12664 29582
rect 12728 22094 12756 32846
rect 12820 31754 12848 33374
rect 12900 32904 12952 32910
rect 12900 32846 12952 32852
rect 12912 32502 12940 32846
rect 13188 32502 13216 33458
rect 12900 32496 12952 32502
rect 12900 32438 12952 32444
rect 13176 32496 13228 32502
rect 13176 32438 13228 32444
rect 13280 32337 13308 35974
rect 13464 35766 13492 37606
rect 13544 37256 13596 37262
rect 13544 37198 13596 37204
rect 13556 36174 13584 37198
rect 13924 36922 13952 39200
rect 14476 37126 14504 39200
rect 14648 37256 14700 37262
rect 14648 37198 14700 37204
rect 14464 37120 14516 37126
rect 14464 37062 14516 37068
rect 13912 36916 13964 36922
rect 13912 36858 13964 36864
rect 14660 36854 14688 37198
rect 15028 37108 15056 39200
rect 15384 37256 15436 37262
rect 15384 37198 15436 37204
rect 15200 37120 15252 37126
rect 15028 37080 15200 37108
rect 15200 37062 15252 37068
rect 14648 36848 14700 36854
rect 14648 36790 14700 36796
rect 14280 36780 14332 36786
rect 14280 36722 14332 36728
rect 14292 36378 14320 36722
rect 14280 36372 14332 36378
rect 14280 36314 14332 36320
rect 15396 36242 15424 37198
rect 15580 36922 15608 39200
rect 15844 37256 15896 37262
rect 15844 37198 15896 37204
rect 15568 36916 15620 36922
rect 15568 36858 15620 36864
rect 15384 36236 15436 36242
rect 15384 36178 15436 36184
rect 13544 36168 13596 36174
rect 13544 36110 13596 36116
rect 15752 36168 15804 36174
rect 15752 36110 15804 36116
rect 13636 36100 13688 36106
rect 13636 36042 13688 36048
rect 13452 35760 13504 35766
rect 13452 35702 13504 35708
rect 13544 35488 13596 35494
rect 13544 35430 13596 35436
rect 13556 34746 13584 35430
rect 13544 34740 13596 34746
rect 13544 34682 13596 34688
rect 13360 33652 13412 33658
rect 13360 33594 13412 33600
rect 13266 32328 13322 32337
rect 13266 32263 13322 32272
rect 13372 31754 13400 33594
rect 13648 31793 13676 36042
rect 13728 35692 13780 35698
rect 13728 35634 13780 35640
rect 13740 34746 13768 35634
rect 14740 35624 14792 35630
rect 14740 35566 14792 35572
rect 14832 35624 14884 35630
rect 14832 35566 14884 35572
rect 14004 35488 14056 35494
rect 14004 35430 14056 35436
rect 13820 35216 13872 35222
rect 13820 35158 13872 35164
rect 13728 34740 13780 34746
rect 13728 34682 13780 34688
rect 13832 33998 13860 35158
rect 14016 35086 14044 35430
rect 14752 35290 14780 35566
rect 14740 35284 14792 35290
rect 14740 35226 14792 35232
rect 14844 35086 14872 35566
rect 15660 35216 15712 35222
rect 15660 35158 15712 35164
rect 15672 35086 15700 35158
rect 14004 35080 14056 35086
rect 14004 35022 14056 35028
rect 14832 35080 14884 35086
rect 14832 35022 14884 35028
rect 15660 35080 15712 35086
rect 15660 35022 15712 35028
rect 14648 34944 14700 34950
rect 14648 34886 14700 34892
rect 14740 34944 14792 34950
rect 14740 34886 14792 34892
rect 14660 34746 14688 34886
rect 14648 34740 14700 34746
rect 14648 34682 14700 34688
rect 14752 34678 14780 34886
rect 15016 34740 15068 34746
rect 15016 34682 15068 34688
rect 14740 34672 14792 34678
rect 14740 34614 14792 34620
rect 14924 34604 14976 34610
rect 14924 34546 14976 34552
rect 14096 34536 14148 34542
rect 14096 34478 14148 34484
rect 14108 33998 14136 34478
rect 14936 34474 14964 34546
rect 14924 34468 14976 34474
rect 14924 34410 14976 34416
rect 14936 34066 14964 34410
rect 14924 34060 14976 34066
rect 14924 34002 14976 34008
rect 13820 33992 13872 33998
rect 13820 33934 13872 33940
rect 14096 33992 14148 33998
rect 14096 33934 14148 33940
rect 13832 33590 13860 33934
rect 13820 33584 13872 33590
rect 13820 33526 13872 33532
rect 14108 33522 14136 33934
rect 15028 33930 15056 34682
rect 15672 34678 15700 35022
rect 15660 34672 15712 34678
rect 15660 34614 15712 34620
rect 15200 34536 15252 34542
rect 15200 34478 15252 34484
rect 15108 34196 15160 34202
rect 15108 34138 15160 34144
rect 15016 33924 15068 33930
rect 15016 33866 15068 33872
rect 14096 33516 14148 33522
rect 14096 33458 14148 33464
rect 15120 33318 15148 34138
rect 15212 33930 15240 34478
rect 15200 33924 15252 33930
rect 15200 33866 15252 33872
rect 14372 33312 14424 33318
rect 14372 33254 14424 33260
rect 15108 33312 15160 33318
rect 15108 33254 15160 33260
rect 14188 32768 14240 32774
rect 14188 32710 14240 32716
rect 14200 32502 14228 32710
rect 14188 32496 14240 32502
rect 14188 32438 14240 32444
rect 13912 32428 13964 32434
rect 13912 32370 13964 32376
rect 13924 32230 13952 32370
rect 13912 32224 13964 32230
rect 13912 32166 13964 32172
rect 13924 32026 13952 32166
rect 13912 32020 13964 32026
rect 13912 31962 13964 31968
rect 13634 31784 13690 31793
rect 12820 31726 12940 31754
rect 13372 31726 13492 31754
rect 12808 30592 12860 30598
rect 12808 30534 12860 30540
rect 12820 30394 12848 30534
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12808 29708 12860 29714
rect 12808 29650 12860 29656
rect 12820 27538 12848 29650
rect 12912 29510 12940 31726
rect 12900 29504 12952 29510
rect 12900 29446 12952 29452
rect 13176 29300 13228 29306
rect 13176 29242 13228 29248
rect 13188 29209 13216 29242
rect 13174 29200 13230 29209
rect 12992 29164 13044 29170
rect 13174 29135 13230 29144
rect 12992 29106 13044 29112
rect 13004 28218 13032 29106
rect 12992 28212 13044 28218
rect 12992 28154 13044 28160
rect 13268 28076 13320 28082
rect 13268 28018 13320 28024
rect 12808 27532 12860 27538
rect 12808 27474 12860 27480
rect 12820 27112 12848 27474
rect 12820 27084 12940 27112
rect 12912 26926 12940 27084
rect 13176 26988 13228 26994
rect 13176 26930 13228 26936
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 12912 26382 12940 26862
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 13188 26314 13216 26930
rect 13176 26308 13228 26314
rect 13176 26250 13228 26256
rect 12728 22066 12940 22094
rect 12268 12406 12388 12434
rect 12544 12406 12664 12434
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11992 9110 12020 9454
rect 11980 9104 12032 9110
rect 11980 9046 12032 9052
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10888 5370 10916 5646
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10520 5273 10548 5306
rect 10506 5264 10562 5273
rect 10980 5234 11008 8774
rect 11992 8430 12020 9046
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 5817 11100 6598
rect 11058 5808 11114 5817
rect 11058 5743 11114 5752
rect 10506 5199 10562 5208
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10428 4282 10456 4558
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10428 3777 10456 4014
rect 10414 3768 10470 3777
rect 10414 3703 10470 3712
rect 10244 3590 10364 3618
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 9954 3224 10010 3233
rect 9954 3159 10010 3168
rect 9968 2922 9996 3159
rect 10060 3058 10088 3334
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 10152 2774 10180 3470
rect 10244 3058 10272 3590
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10060 2746 10180 2774
rect 9954 2680 10010 2689
rect 9954 2615 9956 2624
rect 10008 2615 10010 2624
rect 9956 2586 10008 2592
rect 9864 2100 9916 2106
rect 9864 2042 9916 2048
rect 9310 2000 9366 2009
rect 9310 1935 9366 1944
rect 9496 1760 9548 1766
rect 9496 1702 9548 1708
rect 9508 800 9536 1702
rect 10060 800 10088 2746
rect 10520 2446 10548 4966
rect 10704 4282 10732 5034
rect 10980 5030 11008 5170
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10598 4040 10654 4049
rect 10598 3975 10600 3984
rect 10652 3975 10654 3984
rect 10600 3946 10652 3952
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10704 2774 10732 2994
rect 10888 2990 10916 3334
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10612 2746 10732 2774
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10612 800 10640 2746
rect 10980 2106 11008 4422
rect 11072 2514 11100 5743
rect 11164 3534 11192 7890
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 12084 7546 12112 7754
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11532 6798 11560 7142
rect 11702 7032 11758 7041
rect 11702 6967 11758 6976
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11716 6662 11744 6967
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 12176 6458 12204 7346
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11716 5234 11744 6258
rect 12084 5914 12112 6326
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12176 5030 12204 5170
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11532 3534 11560 4082
rect 11992 3641 12020 4422
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 11978 3632 12034 3641
rect 11704 3596 11756 3602
rect 11978 3567 12034 3576
rect 11704 3538 11756 3544
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11532 3369 11560 3470
rect 11518 3360 11574 3369
rect 11518 3295 11574 3304
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 10968 2100 11020 2106
rect 10968 2042 11020 2048
rect 11164 800 11192 2314
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 1834 11652 2246
rect 11612 1828 11664 1834
rect 11612 1770 11664 1776
rect 11716 800 11744 3538
rect 11888 3460 11940 3466
rect 11888 3402 11940 3408
rect 11900 3126 11928 3402
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11808 2582 11836 2994
rect 11888 2984 11940 2990
rect 11992 2972 12020 3567
rect 11940 2944 12020 2972
rect 11888 2926 11940 2932
rect 12084 2666 12112 4082
rect 12176 3602 12204 4966
rect 12268 4570 12296 12406
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12452 6866 12480 8978
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12360 6254 12388 6734
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12268 4542 12388 4570
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12268 4185 12296 4422
rect 12254 4176 12310 4185
rect 12254 4111 12310 4120
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 12162 3360 12218 3369
rect 12162 3295 12218 3304
rect 11900 2650 12112 2666
rect 11888 2644 12112 2650
rect 11940 2638 12112 2644
rect 11888 2586 11940 2592
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 12176 1442 12204 3295
rect 12268 2582 12296 3878
rect 12360 3777 12388 4542
rect 12452 4146 12480 6802
rect 12544 6390 12572 12406
rect 12808 9512 12860 9518
rect 12806 9480 12808 9489
rect 12860 9480 12862 9489
rect 12806 9415 12862 9424
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12636 8090 12664 8570
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12636 7206 12664 7278
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12636 6730 12664 7142
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 12636 6322 12664 6666
rect 12912 6322 12940 22066
rect 13188 12442 13216 26250
rect 13280 24682 13308 28018
rect 13464 27946 13492 31726
rect 13634 31719 13690 31728
rect 13544 29776 13596 29782
rect 13542 29744 13544 29753
rect 13596 29744 13598 29753
rect 13542 29679 13598 29688
rect 13556 29510 13584 29679
rect 13544 29504 13596 29510
rect 13544 29446 13596 29452
rect 13452 27940 13504 27946
rect 13452 27882 13504 27888
rect 13464 25430 13492 27882
rect 13544 27872 13596 27878
rect 13544 27814 13596 27820
rect 13556 27402 13584 27814
rect 13544 27396 13596 27402
rect 13544 27338 13596 27344
rect 13452 25424 13504 25430
rect 13452 25366 13504 25372
rect 13464 25294 13492 25366
rect 13452 25288 13504 25294
rect 13452 25230 13504 25236
rect 13648 24954 13676 31719
rect 14384 30258 14412 33254
rect 15016 32496 15068 32502
rect 15016 32438 15068 32444
rect 14830 32328 14886 32337
rect 14830 32263 14886 32272
rect 14372 30252 14424 30258
rect 14372 30194 14424 30200
rect 14372 30048 14424 30054
rect 14372 29990 14424 29996
rect 13728 29776 13780 29782
rect 13728 29718 13780 29724
rect 13740 29102 13768 29718
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 14278 29608 14334 29617
rect 13728 29096 13780 29102
rect 13728 29038 13780 29044
rect 14108 28762 14136 29582
rect 14278 29543 14334 29552
rect 14292 29510 14320 29543
rect 14280 29504 14332 29510
rect 14280 29446 14332 29452
rect 14096 28756 14148 28762
rect 14096 28698 14148 28704
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 13820 28416 13872 28422
rect 13820 28358 13872 28364
rect 13832 27538 13860 28358
rect 13820 27532 13872 27538
rect 13820 27474 13872 27480
rect 13832 26330 13860 27474
rect 13740 26302 13860 26330
rect 13740 25498 13768 26302
rect 13820 26240 13872 26246
rect 13820 26182 13872 26188
rect 13728 25492 13780 25498
rect 13728 25434 13780 25440
rect 13636 24948 13688 24954
rect 13636 24890 13688 24896
rect 13452 24744 13504 24750
rect 13452 24686 13504 24692
rect 13268 24676 13320 24682
rect 13268 24618 13320 24624
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13464 11506 13492 24686
rect 13648 24410 13676 24890
rect 13832 24750 13860 26182
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14108 24818 14136 25094
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 13820 24744 13872 24750
rect 13820 24686 13872 24692
rect 14292 24682 14320 28494
rect 14384 26994 14412 29990
rect 14464 27328 14516 27334
rect 14464 27270 14516 27276
rect 14556 27328 14608 27334
rect 14556 27270 14608 27276
rect 14476 27062 14504 27270
rect 14464 27056 14516 27062
rect 14464 26998 14516 27004
rect 14568 26994 14596 27270
rect 14372 26988 14424 26994
rect 14372 26930 14424 26936
rect 14556 26988 14608 26994
rect 14556 26930 14608 26936
rect 14740 26784 14792 26790
rect 14740 26726 14792 26732
rect 14752 26382 14780 26726
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14844 24954 14872 32263
rect 15028 32026 15056 32438
rect 15016 32020 15068 32026
rect 15016 31962 15068 31968
rect 15764 31754 15792 36110
rect 15856 36038 15884 37198
rect 16132 37126 16160 39200
rect 16120 37120 16172 37126
rect 16120 37062 16172 37068
rect 16684 36922 16712 39200
rect 16856 37188 16908 37194
rect 16856 37130 16908 37136
rect 16672 36916 16724 36922
rect 16672 36858 16724 36864
rect 16028 36780 16080 36786
rect 16028 36722 16080 36728
rect 15844 36032 15896 36038
rect 15844 35974 15896 35980
rect 16040 35894 16068 36722
rect 16580 36372 16632 36378
rect 16580 36314 16632 36320
rect 16304 36032 16356 36038
rect 16304 35974 16356 35980
rect 16040 35866 16160 35894
rect 15936 32224 15988 32230
rect 15936 32166 15988 32172
rect 15948 31890 15976 32166
rect 15936 31884 15988 31890
rect 15936 31826 15988 31832
rect 15764 31726 15884 31754
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 15292 30252 15344 30258
rect 15292 30194 15344 30200
rect 15028 28490 15056 30194
rect 15200 30184 15252 30190
rect 15200 30126 15252 30132
rect 15212 29102 15240 30126
rect 15200 29096 15252 29102
rect 15200 29038 15252 29044
rect 15212 28490 15240 29038
rect 15016 28484 15068 28490
rect 15016 28426 15068 28432
rect 15200 28484 15252 28490
rect 15200 28426 15252 28432
rect 15212 28014 15240 28426
rect 15304 28218 15332 30194
rect 15384 29504 15436 29510
rect 15384 29446 15436 29452
rect 15752 29504 15804 29510
rect 15752 29446 15804 29452
rect 15396 29170 15424 29446
rect 15384 29164 15436 29170
rect 15384 29106 15436 29112
rect 15764 29034 15792 29446
rect 15752 29028 15804 29034
rect 15752 28970 15804 28976
rect 15660 28688 15712 28694
rect 15660 28630 15712 28636
rect 15672 28218 15700 28630
rect 15292 28212 15344 28218
rect 15292 28154 15344 28160
rect 15660 28212 15712 28218
rect 15660 28154 15712 28160
rect 15200 28008 15252 28014
rect 15200 27950 15252 27956
rect 14924 27872 14976 27878
rect 14924 27814 14976 27820
rect 14936 27538 14964 27814
rect 15212 27538 15240 27950
rect 14924 27532 14976 27538
rect 14924 27474 14976 27480
rect 15200 27532 15252 27538
rect 15200 27474 15252 27480
rect 14936 26994 14964 27474
rect 15672 27470 15700 28154
rect 15476 27464 15528 27470
rect 15476 27406 15528 27412
rect 15660 27464 15712 27470
rect 15660 27406 15712 27412
rect 15200 27396 15252 27402
rect 15200 27338 15252 27344
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 15212 26790 15240 27338
rect 15200 26784 15252 26790
rect 15200 26726 15252 26732
rect 15488 25498 15516 27406
rect 15568 25696 15620 25702
rect 15568 25638 15620 25644
rect 15476 25492 15528 25498
rect 15476 25434 15528 25440
rect 15016 25356 15068 25362
rect 15016 25298 15068 25304
rect 14832 24948 14884 24954
rect 14832 24890 14884 24896
rect 15028 24750 15056 25298
rect 15580 25226 15608 25638
rect 15568 25220 15620 25226
rect 15568 25162 15620 25168
rect 15292 24812 15344 24818
rect 15292 24754 15344 24760
rect 15016 24744 15068 24750
rect 15016 24686 15068 24692
rect 14280 24676 14332 24682
rect 14280 24618 14332 24624
rect 13636 24404 13688 24410
rect 13636 24346 13688 24352
rect 15304 24070 15332 24754
rect 15292 24064 15344 24070
rect 15292 24006 15344 24012
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13096 11478 13492 11506
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12544 5574 12572 6054
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12452 4010 12480 4082
rect 12440 4004 12492 4010
rect 12440 3946 12492 3952
rect 12346 3768 12402 3777
rect 12346 3703 12402 3712
rect 12544 3512 12572 5510
rect 12636 4826 12664 6258
rect 12898 5944 12954 5953
rect 12898 5879 12900 5888
rect 12952 5879 12954 5888
rect 12992 5908 13044 5914
rect 12900 5850 12952 5856
rect 12992 5850 13044 5856
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12728 4622 12756 5646
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12728 4049 12756 4082
rect 12714 4040 12770 4049
rect 12820 4010 12848 5102
rect 13004 4622 13032 5850
rect 13096 5658 13124 11478
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13372 9450 13400 11086
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13188 5778 13216 6258
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13096 5630 13216 5658
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13004 4282 13032 4558
rect 12992 4276 13044 4282
rect 12992 4218 13044 4224
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 12714 3975 12770 3984
rect 12808 4004 12860 4010
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12532 3506 12584 3512
rect 12532 3448 12584 3454
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12544 3194 12572 3334
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 12360 2310 12388 2586
rect 12636 2446 12664 3606
rect 12728 2774 12756 3975
rect 12808 3946 12860 3952
rect 12820 2990 12848 3946
rect 12912 3534 12940 4150
rect 13004 3602 13032 4218
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 12728 2746 12848 2774
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12452 1902 12480 2382
rect 12440 1896 12492 1902
rect 12440 1838 12492 1844
rect 12636 1766 12664 2382
rect 12624 1760 12676 1766
rect 12624 1702 12676 1708
rect 12176 1414 12296 1442
rect 12268 800 12296 1414
rect 12820 800 12848 2746
rect 13096 1873 13124 4966
rect 13188 4049 13216 5630
rect 13280 4622 13308 8842
rect 13358 6760 13414 6769
rect 13358 6695 13414 6704
rect 13372 6390 13400 6695
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13174 4040 13230 4049
rect 13174 3975 13230 3984
rect 13280 3670 13308 4558
rect 13464 3738 13492 9522
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13556 6322 13584 7346
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13556 5166 13584 6258
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13556 4146 13584 5102
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13542 4040 13598 4049
rect 13542 3975 13598 3984
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13464 2990 13492 3674
rect 13556 3641 13584 3975
rect 13542 3632 13598 3641
rect 13542 3567 13598 3576
rect 13648 3194 13676 11018
rect 13740 9081 13768 12378
rect 14384 11354 14412 13262
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14568 12986 14596 13126
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 15304 12345 15332 24006
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15488 14414 15516 15302
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15672 13938 15700 14214
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15290 12336 15346 12345
rect 15290 12271 15346 12280
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 15198 11248 15254 11257
rect 15198 11183 15254 11192
rect 15212 11150 15240 11183
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 14830 10024 14886 10033
rect 14556 9988 14608 9994
rect 14830 9959 14886 9968
rect 14556 9930 14608 9936
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 13726 9072 13782 9081
rect 13726 9007 13782 9016
rect 13740 8634 13768 9007
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13924 8634 13952 8910
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13740 6322 13768 7346
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14108 6866 14136 7142
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13924 6458 13952 6734
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 14108 5710 14136 6598
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14004 5636 14056 5642
rect 14004 5578 14056 5584
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13740 4593 13768 4694
rect 13726 4584 13782 4593
rect 13726 4519 13782 4528
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13740 3913 13768 4082
rect 13832 4078 13860 5238
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13726 3904 13782 3913
rect 13782 3862 13952 3890
rect 13726 3839 13782 3848
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13648 2854 13676 3130
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 13464 2106 13492 2450
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13556 2106 13584 2246
rect 13452 2100 13504 2106
rect 13452 2042 13504 2048
rect 13544 2100 13596 2106
rect 13544 2042 13596 2048
rect 13740 1902 13768 3334
rect 13832 3058 13860 3334
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13832 2689 13860 2994
rect 13818 2680 13874 2689
rect 13818 2615 13874 2624
rect 13360 1896 13412 1902
rect 13082 1864 13138 1873
rect 13360 1838 13412 1844
rect 13728 1896 13780 1902
rect 13728 1838 13780 1844
rect 13082 1799 13138 1808
rect 13372 800 13400 1838
rect 13924 800 13952 3862
rect 14016 3058 14044 5578
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4622 14228 4966
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14292 4010 14320 8434
rect 14476 7342 14504 9318
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14476 6866 14504 7278
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14384 4622 14412 4966
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14292 3466 14320 3946
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14384 3738 14412 3878
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14476 3534 14504 5578
rect 14568 3602 14596 9930
rect 14844 9110 14872 9959
rect 15304 9654 15332 12271
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15396 11218 15424 11630
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15396 10606 15424 11154
rect 15580 10810 15608 11698
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15764 10742 15792 28970
rect 15856 26042 15884 31726
rect 15936 29708 15988 29714
rect 15936 29650 15988 29656
rect 15948 28014 15976 29650
rect 15936 28008 15988 28014
rect 15936 27950 15988 27956
rect 15844 26036 15896 26042
rect 15844 25978 15896 25984
rect 16132 24342 16160 35866
rect 16212 35692 16264 35698
rect 16212 35634 16264 35640
rect 16224 35222 16252 35634
rect 16212 35216 16264 35222
rect 16212 35158 16264 35164
rect 16316 31906 16344 35974
rect 16488 35488 16540 35494
rect 16488 35430 16540 35436
rect 16500 35222 16528 35430
rect 16488 35216 16540 35222
rect 16488 35158 16540 35164
rect 16396 35148 16448 35154
rect 16396 35090 16448 35096
rect 16408 34134 16436 35090
rect 16396 34128 16448 34134
rect 16396 34070 16448 34076
rect 16500 33930 16528 35158
rect 16592 34406 16620 36314
rect 16868 35894 16896 37130
rect 17236 37126 17264 39200
rect 17788 37330 17816 39200
rect 17776 37324 17828 37330
rect 17776 37266 17828 37272
rect 17684 37256 17736 37262
rect 17684 37198 17736 37204
rect 17224 37120 17276 37126
rect 17224 37062 17276 37068
rect 17696 36825 17724 37198
rect 17682 36816 17738 36825
rect 17040 36780 17092 36786
rect 17682 36751 17738 36760
rect 17040 36722 17092 36728
rect 16776 35866 16896 35894
rect 17052 35894 17080 36722
rect 17696 36310 17724 36751
rect 17788 36378 17816 37266
rect 17972 36802 18000 39222
rect 18248 39114 18276 39222
rect 18326 39200 18382 40000
rect 18878 39200 18934 40000
rect 19430 39200 19486 40000
rect 19982 39200 20038 40000
rect 20534 39200 20590 40000
rect 21086 39200 21142 40000
rect 21638 39200 21694 40000
rect 21744 39222 22048 39250
rect 18340 39114 18368 39200
rect 18248 39086 18368 39114
rect 17880 36786 18000 36802
rect 18604 36848 18656 36854
rect 18604 36790 18656 36796
rect 17868 36780 18000 36786
rect 17920 36774 18000 36780
rect 17868 36722 17920 36728
rect 17868 36576 17920 36582
rect 17868 36518 17920 36524
rect 17776 36372 17828 36378
rect 17776 36314 17828 36320
rect 17684 36304 17736 36310
rect 17684 36246 17736 36252
rect 17052 35866 17448 35894
rect 16672 35624 16724 35630
rect 16672 35566 16724 35572
rect 16684 35222 16712 35566
rect 16672 35216 16724 35222
rect 16672 35158 16724 35164
rect 16580 34400 16632 34406
rect 16580 34342 16632 34348
rect 16684 34202 16712 35158
rect 16776 35086 16804 35866
rect 17236 35834 17264 35866
rect 17224 35828 17276 35834
rect 17224 35770 17276 35776
rect 16764 35080 16816 35086
rect 16764 35022 16816 35028
rect 16672 34196 16724 34202
rect 16672 34138 16724 34144
rect 16776 34082 16804 35022
rect 16856 34400 16908 34406
rect 16856 34342 16908 34348
rect 16592 34054 16804 34082
rect 16592 33930 16620 34054
rect 16488 33924 16540 33930
rect 16488 33866 16540 33872
rect 16580 33924 16632 33930
rect 16580 33866 16632 33872
rect 16500 32230 16528 33866
rect 16592 32298 16620 33866
rect 16672 33856 16724 33862
rect 16672 33798 16724 33804
rect 16684 33522 16712 33798
rect 16672 33516 16724 33522
rect 16672 33458 16724 33464
rect 16764 33312 16816 33318
rect 16764 33254 16816 33260
rect 16776 32434 16804 33254
rect 16764 32428 16816 32434
rect 16764 32370 16816 32376
rect 16580 32292 16632 32298
rect 16580 32234 16632 32240
rect 16488 32224 16540 32230
rect 16488 32166 16540 32172
rect 16316 31878 16436 31906
rect 16304 31816 16356 31822
rect 16304 31758 16356 31764
rect 16316 29306 16344 31758
rect 16304 29300 16356 29306
rect 16304 29242 16356 29248
rect 16212 28416 16264 28422
rect 16212 28358 16264 28364
rect 16224 28082 16252 28358
rect 16212 28076 16264 28082
rect 16212 28018 16264 28024
rect 16120 24336 16172 24342
rect 16120 24278 16172 24284
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 15856 13870 15884 14282
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15948 12850 15976 18022
rect 16224 13433 16252 28018
rect 16408 27033 16436 31878
rect 16672 31340 16724 31346
rect 16672 31282 16724 31288
rect 16684 30326 16712 31282
rect 16868 31113 16896 34342
rect 17040 32292 17092 32298
rect 17040 32234 17092 32240
rect 17052 31278 17080 32234
rect 17132 31884 17184 31890
rect 17132 31826 17184 31832
rect 17040 31272 17092 31278
rect 17040 31214 17092 31220
rect 16854 31104 16910 31113
rect 16854 31039 16910 31048
rect 17144 30802 17172 31826
rect 17132 30796 17184 30802
rect 17132 30738 17184 30744
rect 16672 30320 16724 30326
rect 16486 30288 16542 30297
rect 16672 30262 16724 30268
rect 16486 30223 16542 30232
rect 16500 29850 16528 30223
rect 16488 29844 16540 29850
rect 16488 29786 16540 29792
rect 16500 29646 16528 29786
rect 16488 29640 16540 29646
rect 16488 29582 16540 29588
rect 17224 29504 17276 29510
rect 17224 29446 17276 29452
rect 17236 29306 17264 29446
rect 17224 29300 17276 29306
rect 17224 29242 17276 29248
rect 17224 28552 17276 28558
rect 17224 28494 17276 28500
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 16684 27606 16712 28018
rect 16854 27976 16910 27985
rect 16854 27911 16856 27920
rect 16908 27911 16910 27920
rect 16856 27882 16908 27888
rect 16672 27600 16724 27606
rect 16672 27542 16724 27548
rect 16488 27532 16540 27538
rect 16488 27474 16540 27480
rect 16394 27024 16450 27033
rect 16394 26959 16450 26968
rect 16500 26926 16528 27474
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16488 26920 16540 26926
rect 16488 26862 16540 26868
rect 16396 26784 16448 26790
rect 16396 26726 16448 26732
rect 16304 25220 16356 25226
rect 16304 25162 16356 25168
rect 16210 13424 16266 13433
rect 16210 13359 16266 13368
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 16224 11354 16252 13359
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15396 10130 15424 10542
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 15396 9518 15424 10066
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 14832 9104 14884 9110
rect 14832 9046 14884 9052
rect 14844 8634 14872 9046
rect 15396 8634 15424 9454
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 15120 7857 15148 7958
rect 15200 7880 15252 7886
rect 15106 7848 15162 7857
rect 15200 7822 15252 7828
rect 15106 7783 15162 7792
rect 15212 7546 15240 7822
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15304 7478 15332 8434
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15396 7886 15424 8230
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15488 7528 15516 10610
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15580 8838 15608 10542
rect 15948 10266 15976 11086
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 16316 10033 16344 25162
rect 16408 22030 16436 26726
rect 16500 26382 16528 26862
rect 16960 26790 16988 26930
rect 16948 26784 17000 26790
rect 16948 26726 17000 26732
rect 17144 26586 17172 27406
rect 17132 26580 17184 26586
rect 17132 26522 17184 26528
rect 16488 26376 16540 26382
rect 16488 26318 16540 26324
rect 16948 26376 17000 26382
rect 16948 26318 17000 26324
rect 16960 26042 16988 26318
rect 17132 26308 17184 26314
rect 17132 26250 17184 26256
rect 16948 26036 17000 26042
rect 16948 25978 17000 25984
rect 17040 25968 17092 25974
rect 17038 25936 17040 25945
rect 17092 25936 17094 25945
rect 17038 25871 17094 25880
rect 17144 25838 17172 26250
rect 17132 25832 17184 25838
rect 17132 25774 17184 25780
rect 16488 25764 16540 25770
rect 16488 25706 16540 25712
rect 16500 25362 16528 25706
rect 16670 25664 16726 25673
rect 16670 25599 16726 25608
rect 16488 25356 16540 25362
rect 16488 25298 16540 25304
rect 16684 25294 16712 25599
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 16684 24818 16712 25230
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16948 23656 17000 23662
rect 16948 23598 17000 23604
rect 16960 23322 16988 23598
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 16396 22024 16448 22030
rect 16396 21966 16448 21972
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 16500 17542 16528 18226
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16500 11665 16528 17478
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16592 12238 16620 14214
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16684 12782 16712 13262
rect 16868 12850 16896 16390
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16684 12170 16712 12718
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16486 11656 16542 11665
rect 16408 11614 16486 11642
rect 16302 10024 16358 10033
rect 16302 9959 16358 9968
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15396 7500 15516 7528
rect 15292 7472 15344 7478
rect 15292 7414 15344 7420
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14752 4146 14780 5510
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 14936 4758 14964 5102
rect 15028 5012 15056 5306
rect 15108 5024 15160 5030
rect 15028 4984 15108 5012
rect 15108 4966 15160 4972
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 15120 4690 15148 4966
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 14476 2378 14504 3470
rect 14568 2650 14596 3538
rect 14738 3088 14794 3097
rect 14738 3023 14794 3032
rect 14752 2854 14780 3023
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14844 2650 14872 3538
rect 15108 3460 15160 3466
rect 15108 3402 15160 3408
rect 15120 3194 15148 3402
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 15120 2825 15148 2858
rect 15106 2816 15162 2825
rect 15106 2751 15162 2760
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 15212 2514 15240 4422
rect 15396 4298 15424 7500
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15304 4270 15424 4298
rect 15304 3398 15332 4270
rect 15382 4176 15438 4185
rect 15382 4111 15438 4120
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15396 2990 15424 4111
rect 15488 3942 15516 7346
rect 15580 6866 15608 8774
rect 16408 8634 16436 11614
rect 16486 11591 16542 11600
rect 16592 11150 16620 12038
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16670 11112 16726 11121
rect 16670 11047 16726 11056
rect 16684 10266 16712 11047
rect 16868 10606 16896 12106
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 15948 8498 15976 8570
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 15948 7546 15976 8434
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15948 7342 15976 7482
rect 16500 7342 16528 8502
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 15948 7002 15976 7278
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 16396 6724 16448 6730
rect 16396 6666 16448 6672
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 15750 6216 15806 6225
rect 15750 6151 15806 6160
rect 15764 6118 15792 6151
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15580 5370 15608 6054
rect 15764 5778 15792 6054
rect 16132 5914 16160 6258
rect 16408 6118 16436 6666
rect 16500 6390 16528 7278
rect 16488 6384 16540 6390
rect 16488 6326 16540 6332
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 16408 5234 16436 6054
rect 16500 5778 16528 6326
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 15580 4826 15608 5170
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15672 4622 15700 5170
rect 16488 5160 16540 5166
rect 15842 5128 15898 5137
rect 16488 5102 16540 5108
rect 15842 5063 15898 5072
rect 15856 5030 15884 5063
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 16500 4826 16528 5102
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15936 4548 15988 4554
rect 15936 4490 15988 4496
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 14464 2372 14516 2378
rect 14464 2314 14516 2320
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14200 2038 14228 2246
rect 14188 2032 14240 2038
rect 14188 1974 14240 1980
rect 14464 1760 14516 1766
rect 14464 1702 14516 1708
rect 14476 800 14504 1702
rect 15028 800 15056 2314
rect 15580 800 15608 4082
rect 15672 3670 15700 4218
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 15752 4004 15804 4010
rect 15752 3946 15804 3952
rect 15660 3664 15712 3670
rect 15660 3606 15712 3612
rect 15764 3058 15792 3946
rect 15856 3942 15884 4014
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15948 3194 15976 4490
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16408 3534 16436 4014
rect 16500 3602 16528 4150
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16316 3233 16344 3334
rect 16302 3224 16358 3233
rect 15936 3188 15988 3194
rect 16302 3159 16358 3168
rect 15936 3130 15988 3136
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 16132 800 16160 2790
rect 16592 2106 16620 3674
rect 16684 3466 16712 9862
rect 16960 9217 16988 17274
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 17052 14074 17080 14350
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 17144 12434 17172 25774
rect 17236 24682 17264 28494
rect 17420 26194 17448 35866
rect 17684 33992 17736 33998
rect 17684 33934 17736 33940
rect 17696 33318 17724 33934
rect 17684 33312 17736 33318
rect 17684 33254 17736 33260
rect 17880 32978 17908 36518
rect 17972 35834 18000 36774
rect 18420 36236 18472 36242
rect 18420 36178 18472 36184
rect 17960 35828 18012 35834
rect 17960 35770 18012 35776
rect 18326 33960 18382 33969
rect 18326 33895 18328 33904
rect 18380 33895 18382 33904
rect 18328 33866 18380 33872
rect 18052 33856 18104 33862
rect 18052 33798 18104 33804
rect 18064 33454 18092 33798
rect 18236 33516 18288 33522
rect 18236 33458 18288 33464
rect 18052 33448 18104 33454
rect 18052 33390 18104 33396
rect 18064 33046 18092 33390
rect 18144 33312 18196 33318
rect 18144 33254 18196 33260
rect 18052 33040 18104 33046
rect 18052 32982 18104 32988
rect 17868 32972 17920 32978
rect 17868 32914 17920 32920
rect 17776 31136 17828 31142
rect 17682 31104 17738 31113
rect 17776 31078 17828 31084
rect 17960 31136 18012 31142
rect 17960 31078 18012 31084
rect 17682 31039 17738 31048
rect 17592 30592 17644 30598
rect 17592 30534 17644 30540
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17512 28762 17540 30194
rect 17604 29646 17632 30534
rect 17592 29640 17644 29646
rect 17592 29582 17644 29588
rect 17500 28756 17552 28762
rect 17500 28698 17552 28704
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 17420 26166 17540 26194
rect 17408 25900 17460 25906
rect 17408 25842 17460 25848
rect 17420 25294 17448 25842
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 17512 24954 17540 26166
rect 17500 24948 17552 24954
rect 17500 24890 17552 24896
rect 17500 24744 17552 24750
rect 17500 24686 17552 24692
rect 17224 24676 17276 24682
rect 17224 24618 17276 24624
rect 17512 24070 17540 24686
rect 17500 24064 17552 24070
rect 17500 24006 17552 24012
rect 17408 23316 17460 23322
rect 17408 23258 17460 23264
rect 17420 17218 17448 23258
rect 17512 17338 17540 24006
rect 17604 23866 17632 26930
rect 17696 24886 17724 31039
rect 17788 30938 17816 31078
rect 17776 30932 17828 30938
rect 17776 30874 17828 30880
rect 17972 30734 18000 31078
rect 18064 30870 18092 32982
rect 18156 31142 18184 33254
rect 18248 33114 18276 33458
rect 18236 33108 18288 33114
rect 18236 33050 18288 33056
rect 18144 31136 18196 31142
rect 18144 31078 18196 31084
rect 18052 30864 18104 30870
rect 18052 30806 18104 30812
rect 17960 30728 18012 30734
rect 17960 30670 18012 30676
rect 18052 30660 18104 30666
rect 18052 30602 18104 30608
rect 18064 30054 18092 30602
rect 18052 30048 18104 30054
rect 18052 29990 18104 29996
rect 17868 27328 17920 27334
rect 17868 27270 17920 27276
rect 17880 27062 17908 27270
rect 17868 27056 17920 27062
rect 17868 26998 17920 27004
rect 18144 26988 18196 26994
rect 18144 26930 18196 26936
rect 17960 26784 18012 26790
rect 17960 26726 18012 26732
rect 17972 26450 18000 26726
rect 17960 26444 18012 26450
rect 17960 26386 18012 26392
rect 17960 26240 18012 26246
rect 17960 26182 18012 26188
rect 17972 25838 18000 26182
rect 17960 25832 18012 25838
rect 17960 25774 18012 25780
rect 18156 25362 18184 26930
rect 18328 26784 18380 26790
rect 18328 26726 18380 26732
rect 18340 26314 18368 26726
rect 18328 26308 18380 26314
rect 18328 26250 18380 26256
rect 17960 25356 18012 25362
rect 17960 25298 18012 25304
rect 18144 25356 18196 25362
rect 18144 25298 18196 25304
rect 17684 24880 17736 24886
rect 17684 24822 17736 24828
rect 17696 24410 17724 24822
rect 17972 24750 18000 25298
rect 18052 25152 18104 25158
rect 18052 25094 18104 25100
rect 17960 24744 18012 24750
rect 17960 24686 18012 24692
rect 17684 24404 17736 24410
rect 17684 24346 17736 24352
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17420 17190 17632 17218
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17236 14346 17264 14758
rect 17224 14340 17276 14346
rect 17224 14282 17276 14288
rect 17328 14278 17356 15098
rect 17420 14822 17448 15438
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17420 13870 17448 14758
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17420 13190 17448 13806
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17052 12406 17172 12434
rect 17052 11121 17080 12406
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17038 11112 17094 11121
rect 17038 11047 17094 11056
rect 16946 9208 17002 9217
rect 16946 9143 17002 9152
rect 16960 7546 16988 9143
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16960 7002 16988 7482
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 17052 6322 17080 7686
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16868 5710 16896 6190
rect 16946 5808 17002 5817
rect 16946 5743 17002 5752
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16868 4486 16896 5646
rect 16960 4826 16988 5743
rect 17052 5166 17080 6258
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 17052 4758 17080 5102
rect 17040 4752 17092 4758
rect 17040 4694 17092 4700
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16868 4146 16896 4422
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16776 3534 16804 3878
rect 16868 3602 16896 4082
rect 17144 3738 17172 11698
rect 17236 11150 17264 12582
rect 17328 11150 17356 13126
rect 17512 12374 17540 15370
rect 17500 12368 17552 12374
rect 17500 12310 17552 12316
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17512 11626 17540 12174
rect 17500 11620 17552 11626
rect 17500 11562 17552 11568
rect 17604 11506 17632 17190
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17972 15638 18000 16186
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17788 13326 17816 14214
rect 18064 13462 18092 25094
rect 18340 17241 18368 26250
rect 18432 26042 18460 36178
rect 18616 35894 18644 36790
rect 18892 36174 18920 39200
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 18880 36168 18932 36174
rect 18880 36110 18932 36116
rect 19062 36136 19118 36145
rect 19062 36071 19118 36080
rect 18616 35866 18920 35894
rect 18788 32360 18840 32366
rect 18788 32302 18840 32308
rect 18800 31822 18828 32302
rect 18788 31816 18840 31822
rect 18788 31758 18840 31764
rect 18604 30048 18656 30054
rect 18604 29990 18656 29996
rect 18616 28694 18644 29990
rect 18604 28688 18656 28694
rect 18604 28630 18656 28636
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18524 27130 18552 27406
rect 18512 27124 18564 27130
rect 18512 27066 18564 27072
rect 18512 26512 18564 26518
rect 18512 26454 18564 26460
rect 18420 26036 18472 26042
rect 18420 25978 18472 25984
rect 18432 25537 18460 25978
rect 18418 25528 18474 25537
rect 18418 25463 18474 25472
rect 18432 25294 18460 25463
rect 18420 25288 18472 25294
rect 18420 25230 18472 25236
rect 18524 24206 18552 26454
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18326 17232 18382 17241
rect 18326 17167 18382 17176
rect 18328 17060 18380 17066
rect 18328 17002 18380 17008
rect 18340 16454 18368 17002
rect 18432 16658 18460 17274
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18156 14074 18184 14214
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17788 12782 17816 13126
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17420 11478 17632 11506
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17420 7970 17448 11478
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17512 8974 17540 9318
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17420 7942 17540 7970
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17420 7546 17448 7822
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17406 7440 17462 7449
rect 17406 7375 17462 7384
rect 17420 6662 17448 7375
rect 17512 7206 17540 7942
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17316 6180 17368 6186
rect 17316 6122 17368 6128
rect 17328 5710 17356 6122
rect 17512 5778 17540 7142
rect 17604 5817 17632 11290
rect 17788 9654 17816 12310
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17868 11280 17920 11286
rect 17972 11257 18000 12242
rect 18064 11830 18092 13398
rect 18248 13326 18276 13806
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 18248 12442 18276 13126
rect 18340 12730 18368 16390
rect 18524 13938 18552 16390
rect 18616 16250 18644 28630
rect 18892 28490 18920 35866
rect 19076 30297 19104 36071
rect 19352 35834 19380 37198
rect 19444 36922 19472 39200
rect 19996 37262 20024 39200
rect 20548 37482 20576 39200
rect 20456 37454 20576 37482
rect 20456 37262 20484 37454
rect 21100 37346 21128 39200
rect 21652 39114 21680 39200
rect 21744 39114 21772 39222
rect 21652 39086 21772 39114
rect 21272 37732 21324 37738
rect 21272 37674 21324 37680
rect 21100 37318 21220 37346
rect 21192 37262 21220 37318
rect 19984 37256 20036 37262
rect 19984 37198 20036 37204
rect 20168 37256 20220 37262
rect 20168 37198 20220 37204
rect 20444 37256 20496 37262
rect 20444 37198 20496 37204
rect 21180 37256 21232 37262
rect 21180 37198 21232 37204
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19432 36916 19484 36922
rect 19432 36858 19484 36864
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 19432 36712 19484 36718
rect 19432 36654 19484 36660
rect 19444 36378 19472 36654
rect 19432 36372 19484 36378
rect 19432 36314 19484 36320
rect 19340 35828 19392 35834
rect 19340 35770 19392 35776
rect 19338 35728 19394 35737
rect 19338 35663 19340 35672
rect 19392 35663 19394 35672
rect 19340 35634 19392 35640
rect 19352 35290 19380 35634
rect 19444 35562 19472 36314
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19996 35698 20024 36858
rect 20180 36378 20208 37198
rect 20352 37120 20404 37126
rect 20352 37062 20404 37068
rect 20260 36644 20312 36650
rect 20260 36586 20312 36592
rect 20168 36372 20220 36378
rect 20168 36314 20220 36320
rect 20076 36304 20128 36310
rect 20076 36246 20128 36252
rect 19984 35692 20036 35698
rect 19984 35634 20036 35640
rect 19432 35556 19484 35562
rect 19432 35498 19484 35504
rect 19800 35488 19852 35494
rect 19800 35430 19852 35436
rect 19340 35284 19392 35290
rect 19340 35226 19392 35232
rect 19812 35086 19840 35430
rect 19800 35080 19852 35086
rect 19800 35022 19852 35028
rect 19982 35048 20038 35057
rect 19982 34983 20038 34992
rect 19996 34950 20024 34983
rect 19984 34944 20036 34950
rect 19984 34886 20036 34892
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19432 34536 19484 34542
rect 19432 34478 19484 34484
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19156 32836 19208 32842
rect 19156 32778 19208 32784
rect 19062 30288 19118 30297
rect 19062 30223 19118 30232
rect 18788 28484 18840 28490
rect 18788 28426 18840 28432
rect 18880 28484 18932 28490
rect 18880 28426 18932 28432
rect 18800 28014 18828 28426
rect 18788 28008 18840 28014
rect 18788 27950 18840 27956
rect 18696 27600 18748 27606
rect 18694 27568 18696 27577
rect 18748 27568 18750 27577
rect 18694 27503 18750 27512
rect 18800 26994 18828 27950
rect 18788 26988 18840 26994
rect 18788 26930 18840 26936
rect 18892 24290 18920 28426
rect 18972 28076 19024 28082
rect 18972 28018 19024 28024
rect 18984 25498 19012 28018
rect 19064 26580 19116 26586
rect 19064 26522 19116 26528
rect 19076 26314 19104 26522
rect 19064 26308 19116 26314
rect 19064 26250 19116 26256
rect 19064 26036 19116 26042
rect 19064 25978 19116 25984
rect 19076 25702 19104 25978
rect 19064 25696 19116 25702
rect 19064 25638 19116 25644
rect 18972 25492 19024 25498
rect 18972 25434 19024 25440
rect 19076 24818 19104 25638
rect 19064 24812 19116 24818
rect 19064 24754 19116 24760
rect 18800 24262 18920 24290
rect 18696 24064 18748 24070
rect 18696 24006 18748 24012
rect 18708 23730 18736 24006
rect 18696 23724 18748 23730
rect 18696 23666 18748 23672
rect 18800 23662 18828 24262
rect 18880 24132 18932 24138
rect 18880 24074 18932 24080
rect 18892 23866 18920 24074
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 19076 23526 19104 24754
rect 19064 23520 19116 23526
rect 19064 23462 19116 23468
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18984 16046 19012 16594
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 18984 15570 19012 15982
rect 18972 15564 19024 15570
rect 18972 15506 19024 15512
rect 18984 14958 19012 15506
rect 18972 14952 19024 14958
rect 18892 14900 18972 14906
rect 18892 14894 19024 14900
rect 18892 14878 19012 14894
rect 18892 14482 18920 14878
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 18880 14476 18932 14482
rect 18880 14418 18932 14424
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 18708 13841 18736 14010
rect 18694 13832 18750 13841
rect 18694 13767 18750 13776
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18432 12918 18460 13126
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 18984 12850 19012 14758
rect 19168 14618 19196 32778
rect 19260 27606 19288 32846
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 19352 28218 19380 29106
rect 19340 28212 19392 28218
rect 19340 28154 19392 28160
rect 19248 27600 19300 27606
rect 19248 27542 19300 27548
rect 19260 26382 19288 27542
rect 19340 26920 19392 26926
rect 19340 26862 19392 26868
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19352 23866 19380 26862
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19352 16250 19380 16458
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19444 16182 19472 34478
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 20088 33658 20116 36246
rect 20272 34542 20300 36586
rect 20260 34536 20312 34542
rect 20260 34478 20312 34484
rect 20076 33652 20128 33658
rect 20076 33594 20128 33600
rect 20076 33516 20128 33522
rect 20076 33458 20128 33464
rect 20088 32978 20116 33458
rect 20076 32972 20128 32978
rect 20076 32914 20128 32920
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 20088 31754 20116 32914
rect 20088 31726 20300 31754
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19984 30864 20036 30870
rect 19984 30806 20036 30812
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19996 26586 20024 30806
rect 19616 26580 19668 26586
rect 19616 26522 19668 26528
rect 19984 26580 20036 26586
rect 19984 26522 20036 26528
rect 19522 26480 19578 26489
rect 19522 26415 19524 26424
rect 19576 26415 19578 26424
rect 19524 26386 19576 26392
rect 19628 26246 19656 26522
rect 20168 26444 20220 26450
rect 20168 26386 20220 26392
rect 20076 26308 20128 26314
rect 20076 26250 20128 26256
rect 19616 26240 19668 26246
rect 19616 26182 19668 26188
rect 19984 26240 20036 26246
rect 19984 26182 20036 26188
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19616 24744 19668 24750
rect 19616 24686 19668 24692
rect 19628 24274 19656 24686
rect 19996 24290 20024 26182
rect 20088 25770 20116 26250
rect 20076 25764 20128 25770
rect 20076 25706 20128 25712
rect 20180 25702 20208 26386
rect 20168 25696 20220 25702
rect 20168 25638 20220 25644
rect 20180 25430 20208 25638
rect 20168 25424 20220 25430
rect 20168 25366 20220 25372
rect 20076 25220 20128 25226
rect 20076 25162 20128 25168
rect 20088 24750 20116 25162
rect 20180 24750 20208 25366
rect 20076 24744 20128 24750
rect 20076 24686 20128 24692
rect 20168 24744 20220 24750
rect 20168 24686 20220 24692
rect 19616 24268 19668 24274
rect 19616 24210 19668 24216
rect 19904 24262 20024 24290
rect 20076 24336 20128 24342
rect 20076 24278 20128 24284
rect 19904 24206 19932 24262
rect 19892 24200 19944 24206
rect 19892 24142 19944 24148
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 20088 23866 20116 24278
rect 20076 23860 20128 23866
rect 20076 23802 20128 23808
rect 20088 23769 20116 23802
rect 20074 23760 20130 23769
rect 20074 23695 20130 23704
rect 20180 23662 20208 24686
rect 20168 23656 20220 23662
rect 20168 23598 20220 23604
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 16176 19484 16182
rect 19432 16118 19484 16124
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19168 14278 19196 14554
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19260 13326 19288 15302
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18788 12776 18840 12782
rect 18340 12702 18460 12730
rect 18788 12718 18840 12724
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18156 11898 18184 12174
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18052 11824 18104 11830
rect 18052 11766 18104 11772
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17868 11222 17920 11228
rect 17958 11248 18014 11257
rect 17776 9648 17828 9654
rect 17696 9608 17776 9636
rect 17696 8430 17724 9608
rect 17776 9590 17828 9596
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17788 9382 17816 9454
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 8906 17816 9318
rect 17880 8974 17908 11222
rect 17958 11183 18014 11192
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17776 8900 17828 8906
rect 17776 8842 17828 8848
rect 17960 8560 18012 8566
rect 17960 8502 18012 8508
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17972 7954 18000 8502
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17958 7304 18014 7313
rect 17958 7239 17960 7248
rect 18012 7239 18014 7248
rect 17960 7210 18012 7216
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17788 6118 17816 6190
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17590 5808 17646 5817
rect 17500 5772 17552 5778
rect 17590 5743 17646 5752
rect 17500 5714 17552 5720
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 17236 5302 17264 5510
rect 17224 5296 17276 5302
rect 17224 5238 17276 5244
rect 17236 4146 17264 5238
rect 17328 5098 17356 5646
rect 17512 5642 17540 5714
rect 17500 5636 17552 5642
rect 17500 5578 17552 5584
rect 17960 5636 18012 5642
rect 17960 5578 18012 5584
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17316 5092 17368 5098
rect 17316 5034 17368 5040
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17132 3732 17184 3738
rect 17132 3674 17184 3680
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16684 3097 16712 3402
rect 16670 3088 16726 3097
rect 16670 3023 16726 3032
rect 16868 2990 16896 3538
rect 17420 3194 17448 5170
rect 17972 5166 18000 5578
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 16946 3088 17002 3097
rect 16946 3023 16948 3032
rect 17000 3023 17002 3032
rect 16948 2994 17000 3000
rect 17512 2990 17540 4762
rect 18064 4706 18092 11630
rect 18248 11626 18276 11698
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 18248 10130 18276 11562
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18340 10266 18368 10610
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18432 7528 18460 12702
rect 18800 12442 18828 12718
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18524 11150 18552 12038
rect 19260 11150 19288 12582
rect 19352 12434 19380 14282
rect 19444 12866 19472 15846
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19892 13728 19944 13734
rect 19892 13670 19944 13676
rect 19904 13326 19932 13670
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19444 12838 19564 12866
rect 19996 12850 20024 15302
rect 20088 13818 20116 19654
rect 20180 13938 20208 20198
rect 20272 15162 20300 31726
rect 20364 31414 20392 37062
rect 20456 36106 20484 37198
rect 20812 37188 20864 37194
rect 20812 37130 20864 37136
rect 20824 36922 20852 37130
rect 20904 37120 20956 37126
rect 20904 37062 20956 37068
rect 20996 37120 21048 37126
rect 20996 37062 21048 37068
rect 20812 36916 20864 36922
rect 20812 36858 20864 36864
rect 20628 36236 20680 36242
rect 20628 36178 20680 36184
rect 20444 36100 20496 36106
rect 20444 36042 20496 36048
rect 20444 35692 20496 35698
rect 20444 35634 20496 35640
rect 20456 34678 20484 35634
rect 20640 35222 20668 36178
rect 20628 35216 20680 35222
rect 20628 35158 20680 35164
rect 20640 35086 20668 35158
rect 20628 35080 20680 35086
rect 20628 35022 20680 35028
rect 20720 34944 20772 34950
rect 20720 34886 20772 34892
rect 20732 34678 20760 34886
rect 20444 34672 20496 34678
rect 20444 34614 20496 34620
rect 20720 34672 20772 34678
rect 20720 34614 20772 34620
rect 20444 33992 20496 33998
rect 20444 33934 20496 33940
rect 20456 33658 20484 33934
rect 20444 33652 20496 33658
rect 20444 33594 20496 33600
rect 20732 33538 20760 34614
rect 20916 34474 20944 37062
rect 21008 36854 21036 37062
rect 21284 36938 21312 37674
rect 22020 37210 22048 39222
rect 22190 39200 22246 40000
rect 22742 39200 22798 40000
rect 23294 39200 23350 40000
rect 23846 39200 23902 40000
rect 23952 39222 24256 39250
rect 22112 37262 22140 37293
rect 22100 37256 22152 37262
rect 22020 37204 22100 37210
rect 22020 37198 22152 37204
rect 22020 37182 22140 37198
rect 22204 37194 22232 39200
rect 22112 37074 22140 37182
rect 22192 37188 22244 37194
rect 22192 37130 22244 37136
rect 22112 37046 22232 37074
rect 21192 36922 21312 36938
rect 21180 36916 21312 36922
rect 21232 36910 21312 36916
rect 21180 36858 21232 36864
rect 20996 36848 21048 36854
rect 20996 36790 21048 36796
rect 21192 36553 21220 36858
rect 21548 36712 21600 36718
rect 21548 36654 21600 36660
rect 21178 36544 21234 36553
rect 21178 36479 21234 36488
rect 21086 36408 21142 36417
rect 21086 36343 21142 36352
rect 21100 36038 21128 36343
rect 21560 36242 21588 36654
rect 21730 36272 21786 36281
rect 21548 36236 21600 36242
rect 21730 36207 21786 36216
rect 21548 36178 21600 36184
rect 21272 36100 21324 36106
rect 21272 36042 21324 36048
rect 21088 36032 21140 36038
rect 21088 35974 21140 35980
rect 21100 35834 21128 35974
rect 21088 35828 21140 35834
rect 21088 35770 21140 35776
rect 21088 35488 21140 35494
rect 21088 35430 21140 35436
rect 20904 34468 20956 34474
rect 20904 34410 20956 34416
rect 20640 33510 20760 33538
rect 20640 33454 20668 33510
rect 20628 33448 20680 33454
rect 20628 33390 20680 33396
rect 20732 31890 20760 33510
rect 20812 33312 20864 33318
rect 20812 33254 20864 33260
rect 20824 33153 20852 33254
rect 20810 33144 20866 33153
rect 20810 33079 20866 33088
rect 21100 31890 21128 35430
rect 21284 35086 21312 36042
rect 21560 35630 21588 36178
rect 21744 36106 21772 36207
rect 21732 36100 21784 36106
rect 21732 36042 21784 36048
rect 22100 36100 22152 36106
rect 22100 36042 22152 36048
rect 22112 35834 22140 36042
rect 22100 35828 22152 35834
rect 22100 35770 22152 35776
rect 22204 35714 22232 37046
rect 22374 36544 22430 36553
rect 22374 36479 22430 36488
rect 22388 36174 22416 36479
rect 22376 36168 22428 36174
rect 22376 36110 22428 36116
rect 22560 36168 22612 36174
rect 22560 36110 22612 36116
rect 22572 35834 22600 36110
rect 22756 35873 22784 39200
rect 23308 37346 23336 39200
rect 23860 39114 23888 39200
rect 23952 39114 23980 39222
rect 23860 39086 23980 39114
rect 23848 37732 23900 37738
rect 23848 37674 23900 37680
rect 23860 37466 23888 37674
rect 23848 37460 23900 37466
rect 23848 37402 23900 37408
rect 23308 37318 23428 37346
rect 23296 37256 23348 37262
rect 23296 37198 23348 37204
rect 23112 37120 23164 37126
rect 23112 37062 23164 37068
rect 23020 36712 23072 36718
rect 23020 36654 23072 36660
rect 22742 35864 22798 35873
rect 22560 35828 22612 35834
rect 22742 35799 22798 35808
rect 22560 35770 22612 35776
rect 22112 35686 22232 35714
rect 23032 35714 23060 36654
rect 23124 36242 23152 37062
rect 23112 36236 23164 36242
rect 23112 36178 23164 36184
rect 22744 35692 22796 35698
rect 21548 35624 21600 35630
rect 21548 35566 21600 35572
rect 21638 35184 21694 35193
rect 21638 35119 21694 35128
rect 21272 35080 21324 35086
rect 21272 35022 21324 35028
rect 20720 31884 20772 31890
rect 20720 31826 20772 31832
rect 21088 31884 21140 31890
rect 21088 31826 21140 31832
rect 20732 31754 20760 31826
rect 20732 31726 20852 31754
rect 20352 31408 20404 31414
rect 20352 31350 20404 31356
rect 20444 31340 20496 31346
rect 20444 31282 20496 31288
rect 20456 30938 20484 31282
rect 20824 31278 20852 31726
rect 20720 31272 20772 31278
rect 20720 31214 20772 31220
rect 20812 31272 20864 31278
rect 20812 31214 20864 31220
rect 20444 30932 20496 30938
rect 20444 30874 20496 30880
rect 20732 30734 20760 31214
rect 20536 30728 20588 30734
rect 20536 30670 20588 30676
rect 20720 30728 20772 30734
rect 20772 30688 20852 30716
rect 20720 30670 20772 30676
rect 20548 30326 20576 30670
rect 20536 30320 20588 30326
rect 20536 30262 20588 30268
rect 20534 29336 20590 29345
rect 20534 29271 20590 29280
rect 20548 28626 20576 29271
rect 20824 29238 20852 30688
rect 21088 29640 21140 29646
rect 21088 29582 21140 29588
rect 20996 29572 21048 29578
rect 20996 29514 21048 29520
rect 21008 29481 21036 29514
rect 20994 29472 21050 29481
rect 20994 29407 21050 29416
rect 20812 29232 20864 29238
rect 20812 29174 20864 29180
rect 20996 29232 21048 29238
rect 20996 29174 21048 29180
rect 21008 28914 21036 29174
rect 21100 29102 21128 29582
rect 21088 29096 21140 29102
rect 21088 29038 21140 29044
rect 21180 28960 21232 28966
rect 21008 28886 21128 28914
rect 21180 28902 21232 28908
rect 21100 28626 21128 28886
rect 20536 28620 20588 28626
rect 20536 28562 20588 28568
rect 21088 28620 21140 28626
rect 21088 28562 21140 28568
rect 20548 27878 20576 28562
rect 20536 27872 20588 27878
rect 20536 27814 20588 27820
rect 20548 27334 20576 27814
rect 20812 27464 20864 27470
rect 20812 27406 20864 27412
rect 20720 27396 20772 27402
rect 20720 27338 20772 27344
rect 20536 27328 20588 27334
rect 20536 27270 20588 27276
rect 20548 26994 20576 27270
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 20444 26580 20496 26586
rect 20444 26522 20496 26528
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20364 25430 20392 26318
rect 20352 25424 20404 25430
rect 20352 25366 20404 25372
rect 20352 25152 20404 25158
rect 20352 25094 20404 25100
rect 20364 23254 20392 25094
rect 20456 24857 20484 26522
rect 20548 26042 20576 26930
rect 20626 26480 20682 26489
rect 20626 26415 20682 26424
rect 20536 26036 20588 26042
rect 20536 25978 20588 25984
rect 20536 25764 20588 25770
rect 20536 25706 20588 25712
rect 20442 24848 20498 24857
rect 20442 24783 20498 24792
rect 20352 23248 20404 23254
rect 20352 23190 20404 23196
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 20364 16538 20392 21966
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 20456 19514 20484 19858
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20456 18222 20484 19450
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 20456 16658 20484 18158
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20364 16510 20484 16538
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20364 15162 20392 15438
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20456 15042 20484 16510
rect 20364 15014 20484 15042
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20260 13864 20312 13870
rect 20088 13790 20208 13818
rect 20260 13806 20312 13812
rect 20074 13288 20130 13297
rect 20074 13223 20130 13232
rect 20088 13190 20116 13223
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 19352 12406 19472 12434
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19352 12102 19380 12174
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19352 11082 19380 11562
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18524 9994 18552 10202
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 18512 9988 18564 9994
rect 18512 9930 18564 9936
rect 18604 9988 18656 9994
rect 18604 9930 18656 9936
rect 18524 9722 18552 9930
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 18616 9178 18644 9930
rect 19352 9586 19380 9998
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 18696 9444 18748 9450
rect 18696 9386 18748 9392
rect 18708 9178 18736 9386
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18708 9042 18736 9114
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19352 7970 19380 8978
rect 19168 7954 19380 7970
rect 19168 7948 19392 7954
rect 19168 7942 19340 7948
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18708 7546 18736 7822
rect 18696 7540 18748 7546
rect 18432 7500 18644 7528
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18156 6390 18184 7278
rect 18144 6384 18196 6390
rect 18144 6326 18196 6332
rect 18156 5658 18184 6326
rect 18156 5642 18276 5658
rect 18156 5636 18288 5642
rect 18156 5630 18236 5636
rect 18236 5578 18288 5584
rect 18328 5092 18380 5098
rect 18328 5034 18380 5040
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 17972 4678 18092 4706
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17788 4146 17816 4218
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17604 3194 17632 4082
rect 17972 4078 18000 4678
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 18064 4298 18092 4558
rect 18142 4312 18198 4321
rect 18064 4270 18142 4298
rect 18142 4247 18198 4256
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 18156 3058 18184 4247
rect 18248 4185 18276 4966
rect 18234 4176 18290 4185
rect 18340 4146 18368 5034
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 18234 4111 18290 4120
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 18432 3738 18460 4218
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 16856 2984 16908 2990
rect 16856 2926 16908 2932
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 16580 2100 16632 2106
rect 16580 2042 16632 2048
rect 16684 800 16712 2382
rect 16868 1426 16896 2586
rect 16946 2544 17002 2553
rect 16946 2479 17002 2488
rect 17224 2508 17276 2514
rect 16960 2446 16988 2479
rect 17224 2450 17276 2456
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16960 1834 16988 2382
rect 16948 1828 17000 1834
rect 16948 1770 17000 1776
rect 16856 1420 16908 1426
rect 16856 1362 16908 1368
rect 17236 800 17264 2450
rect 17880 1970 17908 2994
rect 18328 2644 18380 2650
rect 18328 2586 18380 2592
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 17972 2310 18000 2382
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17868 1964 17920 1970
rect 17868 1906 17920 1912
rect 17776 1420 17828 1426
rect 17776 1362 17828 1368
rect 17788 800 17816 1362
rect 18340 800 18368 2586
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18432 2038 18460 2382
rect 18524 2310 18552 7346
rect 18616 7154 18644 7500
rect 18696 7482 18748 7488
rect 18616 7126 18736 7154
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18616 5846 18644 6258
rect 18708 6089 18736 7126
rect 19168 6866 19196 7942
rect 19340 7890 19392 7896
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19260 7002 19288 7822
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 19352 6934 19380 7754
rect 19444 7528 19472 12406
rect 19536 12102 19564 12838
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 19892 12776 19944 12782
rect 19892 12718 19944 12724
rect 19524 12096 19576 12102
rect 19904 12084 19932 12718
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 19904 12056 20024 12084
rect 19524 12038 19576 12044
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19996 10810 20024 12056
rect 19800 10804 19852 10810
rect 19800 10746 19852 10752
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19812 10062 19840 10746
rect 20088 10674 20116 12582
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 20180 10130 20208 13790
rect 20272 12442 20300 13806
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20272 12306 20300 12378
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20168 10124 20220 10130
rect 20168 10066 20220 10072
rect 19800 10056 19852 10062
rect 19800 9998 19852 10004
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 20088 8430 20116 8570
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 20076 8424 20128 8430
rect 20272 8401 20300 10406
rect 20076 8366 20128 8372
rect 20258 8392 20314 8401
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19444 7500 19564 7528
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19340 6928 19392 6934
rect 19340 6870 19392 6876
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 19340 6724 19392 6730
rect 19340 6666 19392 6672
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18984 6458 19012 6598
rect 19352 6458 19380 6666
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19062 6352 19118 6361
rect 19062 6287 19118 6296
rect 18694 6080 18750 6089
rect 18694 6015 18750 6024
rect 18604 5840 18656 5846
rect 18604 5782 18656 5788
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 18616 2854 18644 4626
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 18708 2446 18736 6015
rect 19076 5370 19104 6287
rect 19352 5846 19380 6394
rect 19444 5914 19472 7346
rect 19536 6730 19564 7500
rect 19524 6724 19576 6730
rect 19524 6666 19576 6672
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19340 5840 19392 5846
rect 19168 5788 19340 5794
rect 19168 5782 19392 5788
rect 19168 5766 19380 5782
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18892 3738 18920 5170
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18800 2553 18828 2926
rect 18786 2544 18842 2553
rect 19168 2514 19196 5766
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19352 5234 19380 5578
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19248 4480 19300 4486
rect 19248 4422 19300 4428
rect 19260 3777 19288 4422
rect 19352 4146 19380 5170
rect 19444 4826 19472 5510
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19996 5370 20024 8366
rect 20258 8327 20314 8336
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19246 3768 19302 3777
rect 19246 3703 19302 3712
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19352 3126 19380 3674
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19352 2514 19380 2926
rect 19444 2650 19472 4558
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 19706 3632 19762 3641
rect 19706 3567 19708 3576
rect 19760 3567 19762 3576
rect 19708 3538 19760 3544
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19996 3194 20024 4082
rect 20088 4010 20116 6734
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20180 6458 20208 6598
rect 20168 6452 20220 6458
rect 20168 6394 20220 6400
rect 20260 6180 20312 6186
rect 20260 6122 20312 6128
rect 20272 5642 20300 6122
rect 20260 5636 20312 5642
rect 20260 5578 20312 5584
rect 20272 4826 20300 5578
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20180 4010 20208 4762
rect 20364 4570 20392 15014
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20456 11762 20484 12582
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20548 11642 20576 25706
rect 20640 25294 20668 26415
rect 20628 25288 20680 25294
rect 20628 25230 20680 25236
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20640 24750 20668 25094
rect 20628 24744 20680 24750
rect 20628 24686 20680 24692
rect 20732 24682 20760 27338
rect 20824 27130 20852 27406
rect 20812 27124 20864 27130
rect 20812 27066 20864 27072
rect 20996 25152 21048 25158
rect 20996 25094 21048 25100
rect 21008 24954 21036 25094
rect 20996 24948 21048 24954
rect 20996 24890 21048 24896
rect 20720 24676 20772 24682
rect 20720 24618 20772 24624
rect 20628 23656 20680 23662
rect 20628 23598 20680 23604
rect 20640 23186 20668 23598
rect 20628 23180 20680 23186
rect 20628 23122 20680 23128
rect 20640 22642 20668 23122
rect 20812 23044 20864 23050
rect 20812 22986 20864 22992
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20640 14657 20668 15030
rect 20626 14648 20682 14657
rect 20626 14583 20628 14592
rect 20680 14583 20682 14592
rect 20628 14554 20680 14560
rect 20732 12850 20760 18566
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20628 12708 20680 12714
rect 20628 12650 20680 12656
rect 20640 12209 20668 12650
rect 20626 12200 20682 12209
rect 20626 12135 20682 12144
rect 20548 11614 20668 11642
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 20456 10470 20484 11494
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20548 9042 20576 11494
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20444 8560 20496 8566
rect 20442 8528 20444 8537
rect 20496 8528 20498 8537
rect 20442 8463 20498 8472
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20456 8294 20484 8366
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20456 7954 20484 8230
rect 20444 7948 20496 7954
rect 20444 7890 20496 7896
rect 20456 6186 20484 7890
rect 20444 6180 20496 6186
rect 20444 6122 20496 6128
rect 20536 5840 20588 5846
rect 20536 5782 20588 5788
rect 20548 4622 20576 5782
rect 20536 4616 20588 4622
rect 20364 4542 20484 4570
rect 20536 4558 20588 4564
rect 20076 4004 20128 4010
rect 20076 3946 20128 3952
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 20180 3602 20208 3946
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 20076 3392 20128 3398
rect 20076 3334 20128 3340
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19616 3052 19668 3058
rect 19616 2994 19668 3000
rect 19628 2961 19656 2994
rect 19614 2952 19670 2961
rect 19614 2887 19670 2896
rect 20088 2774 20116 3334
rect 20180 3126 20208 3538
rect 20168 3120 20220 3126
rect 20168 3062 20220 3068
rect 20168 2984 20220 2990
rect 20364 2938 20392 4542
rect 20456 4486 20484 4542
rect 20444 4480 20496 4486
rect 20444 4422 20496 4428
rect 20534 4312 20590 4321
rect 20534 4247 20590 4256
rect 20442 3632 20498 3641
rect 20442 3567 20498 3576
rect 20220 2932 20392 2938
rect 20168 2926 20392 2932
rect 20180 2910 20392 2926
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 19996 2746 20116 2774
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 18786 2479 18842 2488
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 19614 2408 19670 2417
rect 18880 2372 18932 2378
rect 19614 2343 19616 2352
rect 18880 2314 18932 2320
rect 19668 2343 19670 2352
rect 19616 2314 19668 2320
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 18420 2032 18472 2038
rect 18420 1974 18472 1980
rect 18892 800 18920 2314
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19444 800 19472 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2746
rect 20180 2514 20208 2790
rect 20456 2650 20484 3567
rect 20548 3534 20576 4247
rect 20640 3652 20668 11614
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20732 9178 20760 9522
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20824 7834 20852 22986
rect 20996 20800 21048 20806
rect 20996 20742 21048 20748
rect 21008 20602 21036 20742
rect 20996 20596 21048 20602
rect 20996 20538 21048 20544
rect 21100 18426 21128 28562
rect 21192 28558 21220 28902
rect 21180 28552 21232 28558
rect 21180 28494 21232 28500
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 21284 26960 21312 35022
rect 21652 34950 21680 35119
rect 22008 35012 22060 35018
rect 22008 34954 22060 34960
rect 21640 34944 21692 34950
rect 21640 34886 21692 34892
rect 21652 34542 21680 34886
rect 22020 34746 22048 34954
rect 22008 34740 22060 34746
rect 22008 34682 22060 34688
rect 21640 34536 21692 34542
rect 21640 34478 21692 34484
rect 21364 32836 21416 32842
rect 21364 32778 21416 32784
rect 21376 31958 21404 32778
rect 21456 32224 21508 32230
rect 21456 32166 21508 32172
rect 21364 31952 21416 31958
rect 21364 31894 21416 31900
rect 21468 31754 21496 32166
rect 21456 31748 21588 31754
rect 21508 31726 21588 31748
rect 21456 31690 21508 31696
rect 21560 30870 21588 31726
rect 21548 30864 21600 30870
rect 21548 30806 21600 30812
rect 21454 27024 21510 27033
rect 21284 26932 21404 26960
rect 21454 26959 21510 26968
rect 21192 26586 21220 26930
rect 21180 26580 21232 26586
rect 21180 26522 21232 26528
rect 21272 24744 21324 24750
rect 21272 24686 21324 24692
rect 21180 24676 21232 24682
rect 21180 24618 21232 24624
rect 21192 24410 21220 24618
rect 21180 24404 21232 24410
rect 21180 24346 21232 24352
rect 21180 23520 21232 23526
rect 21180 23462 21232 23468
rect 21192 23050 21220 23462
rect 21180 23044 21232 23050
rect 21180 22986 21232 22992
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 21192 19718 21220 19994
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21192 19310 21220 19654
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 21088 18420 21140 18426
rect 21088 18362 21140 18368
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 20916 14890 20944 15302
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 20904 14884 20956 14890
rect 20904 14826 20956 14832
rect 21008 14618 21036 14962
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 21008 14006 21036 14554
rect 20996 14000 21048 14006
rect 20996 13942 21048 13948
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 20916 11694 20944 12786
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20732 7806 20852 7834
rect 20732 7546 20760 7806
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20732 7274 20760 7482
rect 20720 7268 20772 7274
rect 20720 7210 20772 7216
rect 20824 5681 20852 7686
rect 20810 5672 20866 5681
rect 20810 5607 20866 5616
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20732 5370 20760 5510
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20810 4040 20866 4049
rect 20810 3975 20866 3984
rect 20720 3664 20772 3670
rect 20640 3624 20720 3652
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 20076 2372 20128 2378
rect 20076 2314 20128 2320
rect 20088 1902 20116 2314
rect 20076 1896 20128 1902
rect 20076 1838 20128 1844
rect 20548 800 20576 2790
rect 20640 2774 20668 3624
rect 20824 3641 20852 3975
rect 20720 3606 20772 3612
rect 20810 3632 20866 3641
rect 20810 3567 20866 3576
rect 21008 3058 21036 13738
rect 21100 12782 21128 13874
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 21086 9072 21142 9081
rect 21086 9007 21142 9016
rect 21100 8838 21128 9007
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 21100 4826 21128 8366
rect 21088 4820 21140 4826
rect 21088 4762 21140 4768
rect 21100 4214 21128 4762
rect 21088 4208 21140 4214
rect 21088 4150 21140 4156
rect 21192 4146 21220 12718
rect 21284 8430 21312 24686
rect 21376 20058 21404 26932
rect 21468 26382 21496 26959
rect 21456 26376 21508 26382
rect 21456 26318 21508 26324
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21376 19514 21404 19654
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21468 11898 21496 23666
rect 21560 17338 21588 30806
rect 21548 17332 21600 17338
rect 21548 17274 21600 17280
rect 21652 15094 21680 34478
rect 22112 34066 22140 35686
rect 23032 35686 23152 35714
rect 22744 35634 22796 35640
rect 22756 35222 22784 35634
rect 23124 35630 23152 35686
rect 23112 35624 23164 35630
rect 23112 35566 23164 35572
rect 22744 35216 22796 35222
rect 22744 35158 22796 35164
rect 23020 35216 23072 35222
rect 23020 35158 23072 35164
rect 22284 34944 22336 34950
rect 22284 34886 22336 34892
rect 22190 34368 22246 34377
rect 22190 34303 22246 34312
rect 22204 34202 22232 34303
rect 22192 34196 22244 34202
rect 22192 34138 22244 34144
rect 22100 34060 22152 34066
rect 22100 34002 22152 34008
rect 21824 33992 21876 33998
rect 21824 33934 21876 33940
rect 21836 33658 21864 33934
rect 21824 33652 21876 33658
rect 21824 33594 21876 33600
rect 22100 33108 22152 33114
rect 22100 33050 22152 33056
rect 22112 32978 22140 33050
rect 22100 32972 22152 32978
rect 22100 32914 22152 32920
rect 22008 31816 22060 31822
rect 22008 31758 22060 31764
rect 21916 31272 21968 31278
rect 21916 31214 21968 31220
rect 21928 30274 21956 31214
rect 22020 30938 22048 31758
rect 22008 30932 22060 30938
rect 22008 30874 22060 30880
rect 22192 30320 22244 30326
rect 21732 30252 21784 30258
rect 21928 30246 22048 30274
rect 22192 30262 22244 30268
rect 21732 30194 21784 30200
rect 21744 29714 21772 30194
rect 22020 29782 22048 30246
rect 22100 30048 22152 30054
rect 22100 29990 22152 29996
rect 22008 29776 22060 29782
rect 22008 29718 22060 29724
rect 21732 29708 21784 29714
rect 21732 29650 21784 29656
rect 22112 29646 22140 29990
rect 22204 29714 22232 30262
rect 22192 29708 22244 29714
rect 22192 29650 22244 29656
rect 22100 29640 22152 29646
rect 22100 29582 22152 29588
rect 22112 29510 22140 29582
rect 22100 29504 22152 29510
rect 22100 29446 22152 29452
rect 21822 29336 21878 29345
rect 21822 29271 21878 29280
rect 21836 29170 21864 29271
rect 21824 29164 21876 29170
rect 21824 29106 21876 29112
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 21824 28756 21876 28762
rect 21824 28698 21876 28704
rect 21836 28626 21864 28698
rect 21824 28620 21876 28626
rect 21824 28562 21876 28568
rect 21824 27328 21876 27334
rect 21824 27270 21876 27276
rect 21836 27130 21864 27270
rect 21824 27124 21876 27130
rect 21824 27066 21876 27072
rect 21824 25152 21876 25158
rect 21824 25094 21876 25100
rect 21836 24138 21864 25094
rect 21824 24132 21876 24138
rect 21824 24074 21876 24080
rect 21836 23746 21864 24074
rect 21836 23718 21956 23746
rect 21732 22976 21784 22982
rect 21732 22918 21784 22924
rect 21744 22574 21772 22918
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 21732 22568 21784 22574
rect 21732 22510 21784 22516
rect 21836 22030 21864 22578
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 21824 19508 21876 19514
rect 21824 19450 21876 19456
rect 21836 19174 21864 19450
rect 21824 19168 21876 19174
rect 21824 19110 21876 19116
rect 21824 16448 21876 16454
rect 21824 16390 21876 16396
rect 21732 15904 21784 15910
rect 21732 15846 21784 15852
rect 21744 15502 21772 15846
rect 21732 15496 21784 15502
rect 21732 15438 21784 15444
rect 21640 15088 21692 15094
rect 21640 15030 21692 15036
rect 21652 14618 21680 15030
rect 21640 14612 21692 14618
rect 21640 14554 21692 14560
rect 21836 12782 21864 16390
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21652 12345 21680 12378
rect 21638 12336 21694 12345
rect 21638 12271 21694 12280
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21730 11112 21786 11121
rect 21730 11047 21786 11056
rect 21744 11014 21772 11047
rect 21732 11008 21784 11014
rect 21732 10950 21784 10956
rect 21836 10742 21864 12582
rect 21928 11558 21956 23718
rect 22020 23322 22048 29106
rect 22100 26988 22152 26994
rect 22100 26930 22152 26936
rect 22112 24410 22140 26930
rect 22204 26926 22232 29650
rect 22192 26920 22244 26926
rect 22192 26862 22244 26868
rect 22192 26784 22244 26790
rect 22192 26726 22244 26732
rect 22204 26586 22232 26726
rect 22192 26580 22244 26586
rect 22192 26522 22244 26528
rect 22192 25220 22244 25226
rect 22192 25162 22244 25168
rect 22204 24818 22232 25162
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 22100 22568 22152 22574
rect 22100 22510 22152 22516
rect 22112 22030 22140 22510
rect 22296 22094 22324 34886
rect 22560 34604 22612 34610
rect 22560 34546 22612 34552
rect 22572 33658 22600 34546
rect 22560 33652 22612 33658
rect 22560 33594 22612 33600
rect 22742 33552 22798 33561
rect 22742 33487 22744 33496
rect 22796 33487 22798 33496
rect 22928 33516 22980 33522
rect 22744 33458 22796 33464
rect 22928 33458 22980 33464
rect 22756 33046 22784 33458
rect 22744 33040 22796 33046
rect 22742 33008 22744 33017
rect 22796 33008 22798 33017
rect 22742 32943 22798 32952
rect 22742 32872 22798 32881
rect 22742 32807 22798 32816
rect 22468 32428 22520 32434
rect 22468 32370 22520 32376
rect 22480 29170 22508 32370
rect 22756 32298 22784 32807
rect 22744 32292 22796 32298
rect 22744 32234 22796 32240
rect 22560 31136 22612 31142
rect 22560 31078 22612 31084
rect 22572 29646 22600 31078
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22744 29504 22796 29510
rect 22744 29446 22796 29452
rect 22756 29238 22784 29446
rect 22744 29232 22796 29238
rect 22744 29174 22796 29180
rect 22468 29164 22520 29170
rect 22468 29106 22520 29112
rect 22560 27464 22612 27470
rect 22560 27406 22612 27412
rect 22572 27062 22600 27406
rect 22560 27056 22612 27062
rect 22560 26998 22612 27004
rect 22652 27056 22704 27062
rect 22652 26998 22704 27004
rect 22468 26784 22520 26790
rect 22468 26726 22520 26732
rect 22376 26308 22428 26314
rect 22376 26250 22428 26256
rect 22388 24970 22416 26250
rect 22480 25294 22508 26726
rect 22558 25936 22614 25945
rect 22558 25871 22614 25880
rect 22572 25838 22600 25871
rect 22560 25832 22612 25838
rect 22560 25774 22612 25780
rect 22664 25430 22692 26998
rect 22836 26920 22888 26926
rect 22836 26862 22888 26868
rect 22848 26790 22876 26862
rect 22836 26784 22888 26790
rect 22836 26726 22888 26732
rect 22652 25424 22704 25430
rect 22652 25366 22704 25372
rect 22468 25288 22520 25294
rect 22468 25230 22520 25236
rect 22848 25226 22876 26726
rect 22836 25220 22888 25226
rect 22836 25162 22888 25168
rect 22388 24942 22508 24970
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22388 23866 22416 24754
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22480 22094 22508 24942
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22848 23662 22876 24210
rect 22836 23656 22888 23662
rect 22836 23598 22888 23604
rect 22848 23050 22876 23598
rect 22836 23044 22888 23050
rect 22836 22986 22888 22992
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22572 22166 22600 22578
rect 22560 22160 22612 22166
rect 22560 22102 22612 22108
rect 22204 22066 22324 22094
rect 22388 22066 22508 22094
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22112 21010 22140 21830
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 22100 20392 22152 20398
rect 22100 20334 22152 20340
rect 22112 19922 22140 20334
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 22008 19712 22060 19718
rect 22008 19654 22060 19660
rect 22020 16114 22048 19654
rect 22112 19378 22140 19858
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22112 18834 22140 19314
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 22204 15706 22232 22066
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22204 13802 22232 14962
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 22204 13190 22232 13738
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 22388 12434 22416 22066
rect 22940 20058 22968 33458
rect 23032 31754 23060 35158
rect 23124 34082 23152 35566
rect 23204 34604 23256 34610
rect 23204 34546 23256 34552
rect 23216 34202 23244 34546
rect 23204 34196 23256 34202
rect 23204 34138 23256 34144
rect 23124 34066 23244 34082
rect 23124 34060 23256 34066
rect 23124 34054 23204 34060
rect 23204 34002 23256 34008
rect 23112 33856 23164 33862
rect 23112 33798 23164 33804
rect 23124 32774 23152 33798
rect 23216 33454 23244 34002
rect 23204 33448 23256 33454
rect 23204 33390 23256 33396
rect 23308 33046 23336 37198
rect 23400 37194 23428 37318
rect 23664 37256 23716 37262
rect 23664 37198 23716 37204
rect 23388 37188 23440 37194
rect 23388 37130 23440 37136
rect 23676 36922 23704 37198
rect 24122 36952 24178 36961
rect 23664 36916 23716 36922
rect 24122 36887 24178 36896
rect 23664 36858 23716 36864
rect 23386 36816 23442 36825
rect 23386 36751 23388 36760
rect 23440 36751 23442 36760
rect 23388 36722 23440 36728
rect 23480 36712 23532 36718
rect 23386 36680 23442 36689
rect 23480 36654 23532 36660
rect 23386 36615 23388 36624
rect 23440 36615 23442 36624
rect 23388 36586 23440 36592
rect 23492 36242 23520 36654
rect 23756 36576 23808 36582
rect 23756 36518 23808 36524
rect 23768 36310 23796 36518
rect 23756 36304 23808 36310
rect 23756 36246 23808 36252
rect 23480 36236 23532 36242
rect 23480 36178 23532 36184
rect 23388 35692 23440 35698
rect 23388 35634 23440 35640
rect 23400 35465 23428 35634
rect 23386 35456 23442 35465
rect 23386 35391 23442 35400
rect 23400 34950 23428 35391
rect 23664 35284 23716 35290
rect 23664 35226 23716 35232
rect 23388 34944 23440 34950
rect 23388 34886 23440 34892
rect 23386 34776 23442 34785
rect 23386 34711 23388 34720
rect 23440 34711 23442 34720
rect 23388 34682 23440 34688
rect 23676 33386 23704 35226
rect 24136 34513 24164 36887
rect 24228 36854 24256 39222
rect 24398 39200 24454 40000
rect 24950 39200 25006 40000
rect 25502 39200 25558 40000
rect 26054 39200 26110 40000
rect 26606 39200 26662 40000
rect 27158 39200 27214 40000
rect 27710 39200 27766 40000
rect 28262 39200 28318 40000
rect 28814 39200 28870 40000
rect 29366 39200 29422 40000
rect 29918 39200 29974 40000
rect 30470 39200 30526 40000
rect 31022 39200 31078 40000
rect 31128 39222 31432 39250
rect 24216 36848 24268 36854
rect 24216 36790 24268 36796
rect 24412 36258 24440 39200
rect 24676 37120 24728 37126
rect 24676 37062 24728 37068
rect 24688 36961 24716 37062
rect 24674 36952 24730 36961
rect 24674 36887 24730 36896
rect 24768 36848 24820 36854
rect 24768 36790 24820 36796
rect 24412 36230 24532 36258
rect 24400 36168 24452 36174
rect 24400 36110 24452 36116
rect 24306 36000 24362 36009
rect 24306 35935 24362 35944
rect 24320 34746 24348 35935
rect 24412 35834 24440 36110
rect 24400 35828 24452 35834
rect 24400 35770 24452 35776
rect 24504 35086 24532 36230
rect 24582 36136 24638 36145
rect 24582 36071 24638 36080
rect 24596 36038 24624 36071
rect 24584 36032 24636 36038
rect 24584 35974 24636 35980
rect 24492 35080 24544 35086
rect 24492 35022 24544 35028
rect 24492 34944 24544 34950
rect 24492 34886 24544 34892
rect 24308 34740 24360 34746
rect 24308 34682 24360 34688
rect 24122 34504 24178 34513
rect 24122 34439 24178 34448
rect 24032 33856 24084 33862
rect 24032 33798 24084 33804
rect 23664 33380 23716 33386
rect 23664 33322 23716 33328
rect 23296 33040 23348 33046
rect 23296 32982 23348 32988
rect 23112 32768 23164 32774
rect 23112 32710 23164 32716
rect 23386 32600 23442 32609
rect 23386 32535 23442 32544
rect 23400 32502 23428 32535
rect 23388 32496 23440 32502
rect 23388 32438 23440 32444
rect 23032 31726 23336 31754
rect 23112 31680 23164 31686
rect 23112 31622 23164 31628
rect 23124 31414 23152 31622
rect 23112 31408 23164 31414
rect 23112 31350 23164 31356
rect 23204 26784 23256 26790
rect 23204 26726 23256 26732
rect 23020 26308 23072 26314
rect 23020 26250 23072 26256
rect 23032 25974 23060 26250
rect 23020 25968 23072 25974
rect 23020 25910 23072 25916
rect 23216 24614 23244 26726
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 23020 23588 23072 23594
rect 23020 23530 23072 23536
rect 23032 23118 23060 23530
rect 23020 23112 23072 23118
rect 23020 23054 23072 23060
rect 23112 22976 23164 22982
rect 23112 22918 23164 22924
rect 23124 22778 23152 22918
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 23308 20534 23336 31726
rect 23756 26512 23808 26518
rect 23756 26454 23808 26460
rect 23768 25294 23796 26454
rect 23756 25288 23808 25294
rect 23662 25256 23718 25265
rect 23756 25230 23808 25236
rect 23662 25191 23718 25200
rect 23676 25158 23704 25191
rect 23664 25152 23716 25158
rect 23664 25094 23716 25100
rect 23480 24744 23532 24750
rect 23480 24686 23532 24692
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23400 24410 23428 24550
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23388 24268 23440 24274
rect 23388 24210 23440 24216
rect 23400 24070 23428 24210
rect 23388 24064 23440 24070
rect 23388 24006 23440 24012
rect 23492 23730 23520 24686
rect 23572 24608 23624 24614
rect 23572 24550 23624 24556
rect 23584 23866 23612 24550
rect 23676 24138 23704 25094
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23664 24132 23716 24138
rect 23664 24074 23716 24080
rect 23768 23866 23796 24142
rect 23572 23860 23624 23866
rect 23572 23802 23624 23808
rect 23756 23860 23808 23866
rect 23756 23802 23808 23808
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23296 20528 23348 20534
rect 23296 20470 23348 20476
rect 22928 20052 22980 20058
rect 22928 19994 22980 20000
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 23400 16590 23428 18770
rect 23388 16584 23440 16590
rect 23308 16546 23388 16574
rect 22744 16516 22796 16522
rect 22744 16458 22796 16464
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22572 15502 22600 15846
rect 22560 15496 22612 15502
rect 22560 15438 22612 15444
rect 22664 15434 22692 15982
rect 22652 15428 22704 15434
rect 22652 15370 22704 15376
rect 22664 14958 22692 15370
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22664 13938 22692 14894
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22388 12406 22508 12434
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 21916 11552 21968 11558
rect 21916 11494 21968 11500
rect 21824 10736 21876 10742
rect 21824 10678 21876 10684
rect 21822 10024 21878 10033
rect 21822 9959 21878 9968
rect 21836 9926 21864 9959
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21824 9920 21876 9926
rect 21824 9862 21876 9868
rect 21376 9722 21404 9862
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 21560 9110 21588 9454
rect 22204 9450 22232 11698
rect 22480 11558 22508 12406
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22480 10266 22508 11494
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 22192 9444 22244 9450
rect 22192 9386 22244 9392
rect 21548 9104 21600 9110
rect 21548 9046 21600 9052
rect 21732 8900 21784 8906
rect 22756 8888 22784 16458
rect 23308 16046 23336 16546
rect 23388 16526 23440 16532
rect 23296 16040 23348 16046
rect 23296 15982 23348 15988
rect 23308 15570 23336 15982
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23020 13320 23072 13326
rect 23020 13262 23072 13268
rect 22928 13252 22980 13258
rect 22928 13194 22980 13200
rect 22940 12986 22968 13194
rect 22928 12980 22980 12986
rect 22928 12922 22980 12928
rect 23032 12730 23060 13262
rect 23204 12776 23256 12782
rect 23032 12724 23204 12730
rect 23032 12718 23256 12724
rect 23032 12702 23244 12718
rect 23032 12238 23060 12702
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23216 11694 23244 12174
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23204 11688 23256 11694
rect 23400 11665 23428 12038
rect 23204 11630 23256 11636
rect 23386 11656 23442 11665
rect 23216 11150 23244 11630
rect 23386 11591 23442 11600
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 23216 10538 23244 11086
rect 23204 10532 23256 10538
rect 23204 10474 23256 10480
rect 23216 10130 23244 10474
rect 23386 10160 23442 10169
rect 23204 10124 23256 10130
rect 23386 10095 23442 10104
rect 23204 10066 23256 10072
rect 23216 9654 23244 10066
rect 23400 9654 23428 10095
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23492 9602 23520 23666
rect 23584 22094 23612 23802
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 23860 22710 23888 23054
rect 23848 22704 23900 22710
rect 23848 22646 23900 22652
rect 23584 22066 23704 22094
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23584 9926 23612 14758
rect 23676 12646 23704 22066
rect 24044 16182 24072 33798
rect 24136 33289 24164 34439
rect 24504 33658 24532 34886
rect 24582 34096 24638 34105
rect 24780 34066 24808 36790
rect 24860 36032 24912 36038
rect 24860 35974 24912 35980
rect 24872 35494 24900 35974
rect 24860 35488 24912 35494
rect 24860 35430 24912 35436
rect 24964 35086 24992 39200
rect 25136 37256 25188 37262
rect 25320 37256 25372 37262
rect 25188 37204 25320 37210
rect 25136 37198 25372 37204
rect 25148 37182 25360 37198
rect 25044 37120 25096 37126
rect 25044 37062 25096 37068
rect 25136 37120 25188 37126
rect 25136 37062 25188 37068
rect 25320 37120 25372 37126
rect 25320 37062 25372 37068
rect 25056 35766 25084 37062
rect 25148 35873 25176 37062
rect 25332 36242 25360 37062
rect 25412 36916 25464 36922
rect 25412 36858 25464 36864
rect 25424 36689 25452 36858
rect 25516 36802 25544 39200
rect 25778 36816 25834 36825
rect 25516 36774 25728 36802
rect 25504 36712 25556 36718
rect 25410 36680 25466 36689
rect 25504 36654 25556 36660
rect 25410 36615 25466 36624
rect 25320 36236 25372 36242
rect 25320 36178 25372 36184
rect 25516 36174 25544 36654
rect 25504 36168 25556 36174
rect 25504 36110 25556 36116
rect 25228 36032 25280 36038
rect 25228 35974 25280 35980
rect 25134 35864 25190 35873
rect 25134 35799 25190 35808
rect 25044 35760 25096 35766
rect 25044 35702 25096 35708
rect 25240 35222 25268 35974
rect 25516 35698 25544 36110
rect 25700 35698 25728 36774
rect 25778 36751 25834 36760
rect 25320 35692 25372 35698
rect 25320 35634 25372 35640
rect 25504 35692 25556 35698
rect 25504 35634 25556 35640
rect 25688 35692 25740 35698
rect 25688 35634 25740 35640
rect 25332 35290 25360 35634
rect 25410 35456 25466 35465
rect 25410 35391 25466 35400
rect 25320 35284 25372 35290
rect 25320 35226 25372 35232
rect 25424 35222 25452 35391
rect 25228 35216 25280 35222
rect 25228 35158 25280 35164
rect 25412 35216 25464 35222
rect 25412 35158 25464 35164
rect 24952 35080 25004 35086
rect 24952 35022 25004 35028
rect 24860 34604 24912 34610
rect 24860 34546 24912 34552
rect 24582 34031 24584 34040
rect 24636 34031 24638 34040
rect 24768 34060 24820 34066
rect 24584 34002 24636 34008
rect 24768 34002 24820 34008
rect 24596 33862 24624 34002
rect 24584 33856 24636 33862
rect 24584 33798 24636 33804
rect 24492 33652 24544 33658
rect 24492 33594 24544 33600
rect 24122 33280 24178 33289
rect 24122 33215 24178 33224
rect 24400 33040 24452 33046
rect 24400 32982 24452 32988
rect 24412 32842 24440 32982
rect 24400 32836 24452 32842
rect 24400 32778 24452 32784
rect 24492 32836 24544 32842
rect 24492 32778 24544 32784
rect 24400 31952 24452 31958
rect 24400 31894 24452 31900
rect 24412 31793 24440 31894
rect 24398 31784 24454 31793
rect 24398 31719 24454 31728
rect 24400 31340 24452 31346
rect 24400 31282 24452 31288
rect 24308 31136 24360 31142
rect 24308 31078 24360 31084
rect 24412 31090 24440 31282
rect 24504 31210 24532 32778
rect 24676 32224 24728 32230
rect 24676 32166 24728 32172
rect 24492 31204 24544 31210
rect 24492 31146 24544 31152
rect 24320 30870 24348 31078
rect 24412 31062 24532 31090
rect 24308 30864 24360 30870
rect 24308 30806 24360 30812
rect 24400 30048 24452 30054
rect 24400 29990 24452 29996
rect 24412 29850 24440 29990
rect 24400 29844 24452 29850
rect 24400 29786 24452 29792
rect 24400 29504 24452 29510
rect 24398 29472 24400 29481
rect 24452 29472 24454 29481
rect 24398 29407 24454 29416
rect 24504 29034 24532 31062
rect 24688 29753 24716 32166
rect 24872 31906 24900 34546
rect 24964 34202 24992 35022
rect 25136 34944 25188 34950
rect 25136 34886 25188 34892
rect 24952 34196 25004 34202
rect 24952 34138 25004 34144
rect 25148 33998 25176 34886
rect 25516 34626 25544 35634
rect 25516 34610 25636 34626
rect 25516 34604 25648 34610
rect 25516 34598 25596 34604
rect 25596 34546 25648 34552
rect 25412 34196 25464 34202
rect 25412 34138 25464 34144
rect 25136 33992 25188 33998
rect 25136 33934 25188 33940
rect 24780 31890 24900 31906
rect 24768 31884 24900 31890
rect 24820 31878 24900 31884
rect 24964 31878 25176 31906
rect 24768 31826 24820 31832
rect 24964 31822 24992 31878
rect 24952 31816 25004 31822
rect 24952 31758 25004 31764
rect 25044 31816 25096 31822
rect 25044 31758 25096 31764
rect 24674 29744 24730 29753
rect 24674 29679 24730 29688
rect 24860 29572 24912 29578
rect 24860 29514 24912 29520
rect 24492 29028 24544 29034
rect 24492 28970 24544 28976
rect 24308 27328 24360 27334
rect 24308 27270 24360 27276
rect 24400 27328 24452 27334
rect 24400 27270 24452 27276
rect 24320 26450 24348 27270
rect 24308 26444 24360 26450
rect 24308 26386 24360 26392
rect 24412 25401 24440 27270
rect 24398 25392 24454 25401
rect 24398 25327 24454 25336
rect 24400 25220 24452 25226
rect 24400 25162 24452 25168
rect 24412 22982 24440 25162
rect 24400 22976 24452 22982
rect 24400 22918 24452 22924
rect 24412 22710 24440 22918
rect 24400 22704 24452 22710
rect 24400 22646 24452 22652
rect 24504 22094 24532 28970
rect 24872 28121 24900 29514
rect 25056 29209 25084 31758
rect 25148 29850 25176 31878
rect 25136 29844 25188 29850
rect 25136 29786 25188 29792
rect 25042 29200 25098 29209
rect 25042 29135 25098 29144
rect 24858 28112 24914 28121
rect 24858 28047 24914 28056
rect 25044 27872 25096 27878
rect 24964 27832 25044 27860
rect 24858 27432 24914 27441
rect 24858 27367 24860 27376
rect 24912 27367 24914 27376
rect 24860 27338 24912 27344
rect 24964 25906 24992 27832
rect 25044 27814 25096 27820
rect 25044 27328 25096 27334
rect 25044 27270 25096 27276
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 25056 24342 25084 27270
rect 25226 26888 25282 26897
rect 25226 26823 25282 26832
rect 25240 25906 25268 26823
rect 25228 25900 25280 25906
rect 25228 25842 25280 25848
rect 24860 24336 24912 24342
rect 24860 24278 24912 24284
rect 25044 24336 25096 24342
rect 25044 24278 25096 24284
rect 24872 24138 24900 24278
rect 24860 24132 24912 24138
rect 24860 24074 24912 24080
rect 25056 23798 25084 24278
rect 25044 23792 25096 23798
rect 25044 23734 25096 23740
rect 24584 23724 24636 23730
rect 24584 23666 24636 23672
rect 24596 23322 24624 23666
rect 24676 23588 24728 23594
rect 24676 23530 24728 23536
rect 24584 23316 24636 23322
rect 24584 23258 24636 23264
rect 24688 23118 24716 23530
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 25228 23112 25280 23118
rect 25228 23054 25280 23060
rect 25240 22778 25268 23054
rect 25228 22772 25280 22778
rect 25228 22714 25280 22720
rect 24412 22066 24532 22094
rect 24412 16794 24440 22066
rect 25424 18970 25452 34138
rect 25608 33810 25636 34546
rect 25792 34202 25820 36751
rect 25964 36576 26016 36582
rect 25964 36518 26016 36524
rect 25976 36106 26004 36518
rect 25964 36100 26016 36106
rect 25964 36042 26016 36048
rect 26068 35766 26096 39200
rect 26240 37664 26292 37670
rect 26240 37606 26292 37612
rect 26146 36544 26202 36553
rect 26146 36479 26202 36488
rect 26056 35760 26108 35766
rect 26056 35702 26108 35708
rect 26056 35488 26108 35494
rect 26056 35430 26108 35436
rect 25780 34196 25832 34202
rect 25780 34138 25832 34144
rect 25608 33782 25820 33810
rect 25792 32910 25820 33782
rect 26068 33590 26096 35430
rect 26160 35290 26188 36479
rect 26252 36106 26280 37606
rect 26330 36816 26386 36825
rect 26330 36751 26386 36760
rect 26344 36650 26372 36751
rect 26332 36644 26384 36650
rect 26332 36586 26384 36592
rect 26240 36100 26292 36106
rect 26240 36042 26292 36048
rect 26238 35864 26294 35873
rect 26238 35799 26294 35808
rect 26148 35284 26200 35290
rect 26148 35226 26200 35232
rect 26252 34746 26280 35799
rect 26620 35086 26648 39200
rect 27172 37126 27200 39200
rect 27436 37256 27488 37262
rect 27436 37198 27488 37204
rect 27160 37120 27212 37126
rect 27160 37062 27212 37068
rect 26976 36576 27028 36582
rect 26976 36518 27028 36524
rect 26988 36281 27016 36518
rect 27448 36378 27476 37198
rect 27724 37126 27752 39200
rect 28080 37256 28132 37262
rect 28080 37198 28132 37204
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 27436 36372 27488 36378
rect 27436 36314 27488 36320
rect 26974 36272 27030 36281
rect 26974 36207 27030 36216
rect 27712 36032 27764 36038
rect 27712 35974 27764 35980
rect 27620 35488 27672 35494
rect 27620 35430 27672 35436
rect 26608 35080 26660 35086
rect 26608 35022 26660 35028
rect 26240 34740 26292 34746
rect 26240 34682 26292 34688
rect 26976 34740 27028 34746
rect 26976 34682 27028 34688
rect 26988 34649 27016 34682
rect 26974 34640 27030 34649
rect 26974 34575 27030 34584
rect 26056 33584 26108 33590
rect 26056 33526 26108 33532
rect 27632 33522 27660 35430
rect 27724 35222 27752 35974
rect 27896 35692 27948 35698
rect 27896 35634 27948 35640
rect 27988 35692 28040 35698
rect 27988 35634 28040 35640
rect 27908 35290 27936 35634
rect 27896 35284 27948 35290
rect 27896 35226 27948 35232
rect 27712 35216 27764 35222
rect 27712 35158 27764 35164
rect 28000 34678 28028 35634
rect 28092 34932 28120 37198
rect 28276 37126 28304 39200
rect 28448 37460 28500 37466
rect 28448 37402 28500 37408
rect 28264 37120 28316 37126
rect 28264 37062 28316 37068
rect 28170 36952 28226 36961
rect 28170 36887 28172 36896
rect 28224 36887 28226 36896
rect 28172 36858 28224 36864
rect 28460 36650 28488 37402
rect 28828 37210 28856 39200
rect 29380 37466 29408 39200
rect 29368 37460 29420 37466
rect 29368 37402 29420 37408
rect 29276 37256 29328 37262
rect 28828 37182 29040 37210
rect 29276 37198 29328 37204
rect 29012 37126 29040 37182
rect 29000 37120 29052 37126
rect 29000 37062 29052 37068
rect 29000 36712 29052 36718
rect 29000 36654 29052 36660
rect 28448 36644 28500 36650
rect 28448 36586 28500 36592
rect 29012 36174 29040 36654
rect 29288 36582 29316 37198
rect 29932 37126 29960 39200
rect 30380 37256 30432 37262
rect 30380 37198 30432 37204
rect 30104 37188 30156 37194
rect 30104 37130 30156 37136
rect 29920 37120 29972 37126
rect 29920 37062 29972 37068
rect 29276 36576 29328 36582
rect 29276 36518 29328 36524
rect 29000 36168 29052 36174
rect 29000 36110 29052 36116
rect 28998 35320 29054 35329
rect 28998 35255 29054 35264
rect 28172 34944 28224 34950
rect 28092 34904 28172 34932
rect 28172 34886 28224 34892
rect 27988 34672 28040 34678
rect 27988 34614 28040 34620
rect 28080 34604 28132 34610
rect 28080 34546 28132 34552
rect 27802 34232 27858 34241
rect 27802 34167 27858 34176
rect 27816 33998 27844 34167
rect 27804 33992 27856 33998
rect 27804 33934 27856 33940
rect 27620 33516 27672 33522
rect 27620 33458 27672 33464
rect 27804 33516 27856 33522
rect 27804 33458 27856 33464
rect 26330 33280 26386 33289
rect 26330 33215 26386 33224
rect 25780 32904 25832 32910
rect 25780 32846 25832 32852
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 26068 32434 26096 32846
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 26148 32428 26200 32434
rect 26148 32370 26200 32376
rect 26068 31890 26096 32370
rect 26160 32026 26188 32370
rect 26148 32020 26200 32026
rect 26148 31962 26200 31968
rect 26056 31884 26108 31890
rect 26056 31826 26108 31832
rect 25596 31408 25648 31414
rect 25596 31350 25648 31356
rect 25608 30054 25636 31350
rect 26068 31346 26096 31826
rect 26056 31340 26108 31346
rect 26056 31282 26108 31288
rect 26068 30802 26096 31282
rect 26056 30796 26108 30802
rect 26056 30738 26108 30744
rect 26344 30122 26372 33215
rect 27252 32836 27304 32842
rect 27252 32778 27304 32784
rect 27264 32609 27292 32778
rect 27250 32600 27306 32609
rect 27250 32535 27306 32544
rect 27620 32224 27672 32230
rect 27620 32166 27672 32172
rect 27632 31482 27660 32166
rect 27620 31476 27672 31482
rect 27620 31418 27672 31424
rect 27816 30734 27844 33458
rect 28092 31142 28120 34546
rect 28080 31136 28132 31142
rect 28080 31078 28132 31084
rect 27804 30728 27856 30734
rect 27804 30670 27856 30676
rect 27620 30252 27672 30258
rect 27620 30194 27672 30200
rect 26516 30184 26568 30190
rect 26516 30126 26568 30132
rect 25872 30116 25924 30122
rect 25872 30058 25924 30064
rect 26332 30116 26384 30122
rect 26332 30058 26384 30064
rect 25596 30048 25648 30054
rect 25596 29990 25648 29996
rect 25596 29300 25648 29306
rect 25596 29242 25648 29248
rect 25608 28490 25636 29242
rect 25596 28484 25648 28490
rect 25596 28426 25648 28432
rect 25504 24064 25556 24070
rect 25504 24006 25556 24012
rect 25516 22098 25544 24006
rect 25884 23186 25912 30058
rect 26424 30048 26476 30054
rect 26424 29990 26476 29996
rect 25964 29844 26016 29850
rect 25964 29786 26016 29792
rect 25976 23798 26004 29786
rect 26240 28008 26292 28014
rect 26240 27950 26292 27956
rect 26252 27470 26280 27950
rect 26436 27538 26464 29990
rect 26528 29646 26556 30126
rect 26516 29640 26568 29646
rect 26516 29582 26568 29588
rect 26528 29102 26556 29582
rect 26516 29096 26568 29102
rect 27632 29073 27660 30194
rect 26516 29038 26568 29044
rect 27618 29064 27674 29073
rect 26528 28558 26556 29038
rect 27618 28999 27674 29008
rect 26516 28552 26568 28558
rect 26516 28494 26568 28500
rect 26974 28520 27030 28529
rect 26528 28014 26556 28494
rect 26974 28455 27030 28464
rect 26516 28008 26568 28014
rect 26516 27950 26568 27956
rect 26424 27532 26476 27538
rect 26424 27474 26476 27480
rect 26240 27464 26292 27470
rect 26240 27406 26292 27412
rect 26252 26926 26280 27406
rect 26424 27396 26476 27402
rect 26424 27338 26476 27344
rect 26240 26920 26292 26926
rect 26240 26862 26292 26868
rect 26252 26314 26280 26862
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26252 25838 26280 26250
rect 26240 25832 26292 25838
rect 26240 25774 26292 25780
rect 26252 25294 26280 25774
rect 26240 25288 26292 25294
rect 26240 25230 26292 25236
rect 26332 25220 26384 25226
rect 26332 25162 26384 25168
rect 26344 24274 26372 25162
rect 26436 24410 26464 27338
rect 26988 26858 27016 28455
rect 27620 26988 27672 26994
rect 27620 26930 27672 26936
rect 26976 26852 27028 26858
rect 26976 26794 27028 26800
rect 27632 26353 27660 26930
rect 27816 26382 27844 30670
rect 28184 29510 28212 34886
rect 29012 34202 29040 35255
rect 29092 35148 29144 35154
rect 29092 35090 29144 35096
rect 29104 34746 29132 35090
rect 29092 34740 29144 34746
rect 29092 34682 29144 34688
rect 29184 34740 29236 34746
rect 29184 34682 29236 34688
rect 29196 34377 29224 34682
rect 29182 34368 29238 34377
rect 29182 34303 29238 34312
rect 29000 34196 29052 34202
rect 29000 34138 29052 34144
rect 28998 33144 29054 33153
rect 28998 33079 29054 33088
rect 29012 32910 29040 33079
rect 29000 32904 29052 32910
rect 29000 32846 29052 32852
rect 29288 31754 29316 36518
rect 29460 36236 29512 36242
rect 29460 36178 29512 36184
rect 29288 31726 29408 31754
rect 29000 31340 29052 31346
rect 29000 31282 29052 31288
rect 28356 31136 28408 31142
rect 28354 31104 28356 31113
rect 28408 31104 28410 31113
rect 28354 31039 28410 31048
rect 29012 30326 29040 31282
rect 29092 31136 29144 31142
rect 29092 31078 29144 31084
rect 29000 30320 29052 30326
rect 29000 30262 29052 30268
rect 28356 30252 28408 30258
rect 28356 30194 28408 30200
rect 28172 29504 28224 29510
rect 28172 29446 28224 29452
rect 27988 29028 28040 29034
rect 27988 28970 28040 28976
rect 27804 26376 27856 26382
rect 27618 26344 27674 26353
rect 27804 26318 27856 26324
rect 27618 26279 27674 26288
rect 28000 25537 28028 28970
rect 27986 25528 28042 25537
rect 27986 25463 28042 25472
rect 27710 24848 27766 24857
rect 27710 24783 27766 24792
rect 27724 24682 27752 24783
rect 27712 24676 27764 24682
rect 27712 24618 27764 24624
rect 26424 24404 26476 24410
rect 26424 24346 26476 24352
rect 26332 24268 26384 24274
rect 26332 24210 26384 24216
rect 28080 24200 28132 24206
rect 28080 24142 28132 24148
rect 26148 24064 26200 24070
rect 26148 24006 26200 24012
rect 25964 23792 26016 23798
rect 25964 23734 26016 23740
rect 26160 23662 26188 24006
rect 26608 23792 26660 23798
rect 26608 23734 26660 23740
rect 26056 23656 26108 23662
rect 26056 23598 26108 23604
rect 26148 23656 26200 23662
rect 26148 23598 26200 23604
rect 25872 23180 25924 23186
rect 25872 23122 25924 23128
rect 25596 22636 25648 22642
rect 25596 22578 25648 22584
rect 25608 22234 25636 22578
rect 25596 22228 25648 22234
rect 25596 22170 25648 22176
rect 25504 22092 25556 22098
rect 25504 22034 25556 22040
rect 25412 18964 25464 18970
rect 25412 18906 25464 18912
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 25148 16590 25176 17070
rect 25136 16584 25188 16590
rect 26068 16574 26096 23598
rect 26620 23322 26648 23734
rect 26608 23316 26660 23322
rect 26608 23258 26660 23264
rect 27712 22976 27764 22982
rect 27712 22918 27764 22924
rect 27724 22642 27752 22918
rect 27712 22636 27764 22642
rect 27712 22578 27764 22584
rect 27620 22568 27672 22574
rect 27620 22510 27672 22516
rect 27632 22098 27660 22510
rect 26792 22092 26844 22098
rect 26792 22034 26844 22040
rect 27620 22092 27672 22098
rect 27620 22034 27672 22040
rect 26804 21486 26832 22034
rect 26976 22024 27028 22030
rect 26976 21966 27028 21972
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 26792 21480 26844 21486
rect 26792 21422 26844 21428
rect 26240 18692 26292 18698
rect 26240 18634 26292 18640
rect 26252 16574 26280 18634
rect 26424 17060 26476 17066
rect 26424 17002 26476 17008
rect 26068 16546 26188 16574
rect 26252 16546 26372 16574
rect 25136 16526 25188 16532
rect 24032 16176 24084 16182
rect 24032 16118 24084 16124
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24412 15162 24440 15438
rect 24400 15156 24452 15162
rect 24400 15098 24452 15104
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23768 13802 23796 14010
rect 23756 13796 23808 13802
rect 23756 13738 23808 13744
rect 24492 13456 24544 13462
rect 24490 13424 24492 13433
rect 24544 13424 24546 13433
rect 24490 13359 24546 13368
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 23572 9920 23624 9926
rect 23572 9862 23624 9868
rect 23216 9042 23244 9590
rect 23492 9574 23612 9602
rect 23584 9450 23612 9574
rect 23572 9444 23624 9450
rect 23572 9386 23624 9392
rect 23204 9036 23256 9042
rect 23204 8978 23256 8984
rect 22836 8900 22888 8906
rect 22756 8860 22836 8888
rect 21732 8842 21784 8848
rect 22836 8842 22888 8848
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 21744 8362 21772 8842
rect 22008 8560 22060 8566
rect 22008 8502 22060 8508
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 22020 8294 22048 8502
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22008 8288 22060 8294
rect 22008 8230 22060 8236
rect 22006 7848 22062 7857
rect 22006 7783 22062 7792
rect 22284 7812 22336 7818
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21638 6760 21694 6769
rect 21638 6695 21694 6704
rect 21652 6662 21680 6695
rect 21744 6662 21772 6802
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 22020 6610 22048 7783
rect 22284 7754 22336 7760
rect 22296 7313 22324 7754
rect 22282 7304 22338 7313
rect 22282 7239 22338 7248
rect 22388 7154 22416 8434
rect 22296 7126 22416 7154
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22204 6610 22232 6734
rect 22296 6730 22324 7126
rect 22374 6896 22430 6905
rect 22374 6831 22430 6840
rect 22284 6724 22336 6730
rect 22284 6666 22336 6672
rect 22020 6582 22232 6610
rect 22388 6458 22416 6831
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 21456 6180 21508 6186
rect 21456 6122 21508 6128
rect 21468 5710 21496 6122
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21284 5302 21312 5646
rect 21272 5296 21324 5302
rect 21836 5273 21864 6054
rect 22296 5642 22324 6394
rect 22650 5944 22706 5953
rect 22650 5879 22706 5888
rect 22664 5710 22692 5879
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 22284 5636 22336 5642
rect 22284 5578 22336 5584
rect 21916 5296 21968 5302
rect 21272 5238 21324 5244
rect 21822 5264 21878 5273
rect 21284 4826 21312 5238
rect 21916 5238 21968 5244
rect 21822 5199 21878 5208
rect 21824 5024 21876 5030
rect 21928 5012 21956 5238
rect 21876 4984 21956 5012
rect 21824 4966 21876 4972
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 21640 4480 21692 4486
rect 21640 4422 21692 4428
rect 21284 4146 21312 4422
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 21272 4140 21324 4146
rect 21272 4082 21324 4088
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 21100 3602 21128 3878
rect 21088 3596 21140 3602
rect 21088 3538 21140 3544
rect 21192 3534 21220 4082
rect 21272 3936 21324 3942
rect 21652 3913 21680 4422
rect 21836 4010 21864 4966
rect 22374 4584 22430 4593
rect 22374 4519 22376 4528
rect 22428 4519 22430 4528
rect 22376 4490 22428 4496
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 21824 4004 21876 4010
rect 21824 3946 21876 3952
rect 21272 3878 21324 3884
rect 21638 3904 21694 3913
rect 21284 3670 21312 3878
rect 21638 3839 21694 3848
rect 21272 3664 21324 3670
rect 21272 3606 21324 3612
rect 21180 3528 21232 3534
rect 21180 3470 21232 3476
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21376 3058 21404 3470
rect 22112 3058 22140 4422
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 20996 3052 21048 3058
rect 20996 2994 21048 3000
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 22192 2848 22244 2854
rect 22192 2790 22244 2796
rect 20640 2746 20760 2774
rect 20732 2446 20760 2746
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 21088 2304 21140 2310
rect 21088 2246 21140 2252
rect 21100 800 21128 2246
rect 21640 2100 21692 2106
rect 21640 2042 21692 2048
rect 21652 800 21680 2042
rect 22204 800 22232 2790
rect 22480 2446 22508 3878
rect 22756 3738 22784 4082
rect 22848 3942 22876 8842
rect 23216 8498 23244 8978
rect 23584 8838 23612 9386
rect 23572 8832 23624 8838
rect 23572 8774 23624 8780
rect 23204 8492 23256 8498
rect 23204 8434 23256 8440
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23492 7342 23520 7822
rect 23480 7336 23532 7342
rect 23480 7278 23532 7284
rect 23492 6798 23520 7278
rect 23570 7032 23626 7041
rect 23570 6967 23626 6976
rect 23584 6798 23612 6967
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23492 6254 23520 6734
rect 23480 6248 23532 6254
rect 23480 6190 23532 6196
rect 23492 5710 23520 6190
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 23492 5166 23520 5646
rect 23676 5642 23704 12582
rect 23768 7750 23796 12786
rect 24872 12434 24900 16050
rect 24950 15192 25006 15201
rect 24950 15127 24952 15136
rect 25004 15127 25006 15136
rect 24952 15098 25004 15104
rect 24964 14550 24992 15098
rect 25148 14958 25176 16526
rect 25596 15632 25648 15638
rect 25596 15574 25648 15580
rect 25412 15360 25464 15366
rect 25412 15302 25464 15308
rect 25504 15360 25556 15366
rect 25504 15302 25556 15308
rect 25424 15094 25452 15302
rect 25412 15088 25464 15094
rect 25412 15030 25464 15036
rect 25320 15020 25372 15026
rect 25320 14962 25372 14968
rect 25136 14952 25188 14958
rect 25136 14894 25188 14900
rect 24952 14544 25004 14550
rect 24952 14486 25004 14492
rect 25148 14482 25176 14894
rect 25332 14618 25360 14962
rect 25320 14612 25372 14618
rect 25320 14554 25372 14560
rect 25424 14482 25452 15030
rect 25516 14958 25544 15302
rect 25504 14952 25556 14958
rect 25504 14894 25556 14900
rect 25136 14476 25188 14482
rect 25136 14418 25188 14424
rect 25412 14476 25464 14482
rect 25412 14418 25464 14424
rect 25412 14272 25464 14278
rect 25412 14214 25464 14220
rect 25424 14074 25452 14214
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25424 13938 25452 14010
rect 25412 13932 25464 13938
rect 25412 13874 25464 13880
rect 25516 13870 25544 14010
rect 25504 13864 25556 13870
rect 25504 13806 25556 13812
rect 25504 12844 25556 12850
rect 25504 12786 25556 12792
rect 24872 12406 24992 12434
rect 24768 11076 24820 11082
rect 24768 11018 24820 11024
rect 23848 9920 23900 9926
rect 23848 9862 23900 9868
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 23664 5636 23716 5642
rect 23664 5578 23716 5584
rect 23480 5160 23532 5166
rect 23480 5102 23532 5108
rect 23492 4622 23520 5102
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23492 4146 23520 4558
rect 23584 4282 23612 4558
rect 23860 4554 23888 9862
rect 24780 9382 24808 11018
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 24768 9376 24820 9382
rect 24964 9353 24992 12406
rect 25228 12164 25280 12170
rect 25228 12106 25280 12112
rect 25240 11830 25268 12106
rect 25228 11824 25280 11830
rect 25228 11766 25280 11772
rect 25516 11762 25544 12786
rect 25608 11898 25636 15574
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 26068 14958 26096 15438
rect 26056 14952 26108 14958
rect 26056 14894 26108 14900
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25884 12850 25912 13262
rect 25872 12844 25924 12850
rect 25872 12786 25924 12792
rect 25596 11892 25648 11898
rect 25596 11834 25648 11840
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 25228 11008 25280 11014
rect 25228 10950 25280 10956
rect 25240 9489 25268 10950
rect 25516 10538 25544 11698
rect 26056 10668 26108 10674
rect 26056 10610 26108 10616
rect 25504 10532 25556 10538
rect 25504 10474 25556 10480
rect 25516 9586 25544 10474
rect 26068 10062 26096 10610
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 25504 9580 25556 9586
rect 25504 9522 25556 9528
rect 25226 9480 25282 9489
rect 25226 9415 25282 9424
rect 24768 9318 24820 9324
rect 24950 9344 25006 9353
rect 24044 8945 24072 9318
rect 24950 9279 25006 9288
rect 24030 8936 24086 8945
rect 24030 8871 24086 8880
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 24872 8090 24900 8842
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 24768 6724 24820 6730
rect 24768 6666 24820 6672
rect 24780 6118 24808 6666
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24860 6112 24912 6118
rect 24860 6054 24912 6060
rect 24872 5234 24900 6054
rect 24964 5302 24992 9279
rect 25516 8906 25544 9522
rect 25504 8900 25556 8906
rect 25504 8842 25556 8848
rect 26160 8362 26188 16546
rect 26344 12434 26372 16546
rect 26436 15638 26464 17002
rect 26988 16574 27016 21966
rect 27252 21956 27304 21962
rect 27252 21898 27304 21904
rect 27160 21888 27212 21894
rect 27160 21830 27212 21836
rect 27172 21350 27200 21830
rect 27160 21344 27212 21350
rect 27160 21286 27212 21292
rect 27068 20596 27120 20602
rect 27068 20538 27120 20544
rect 26896 16546 27016 16574
rect 27080 16574 27108 20538
rect 27172 19310 27200 21286
rect 27264 21146 27292 21898
rect 28000 21146 28028 21966
rect 28092 21894 28120 24142
rect 28184 22166 28212 29446
rect 28368 23866 28396 30194
rect 28908 29776 28960 29782
rect 28908 29718 28960 29724
rect 28920 25945 28948 29718
rect 29104 29578 29132 31078
rect 29276 30048 29328 30054
rect 29276 29990 29328 29996
rect 29092 29572 29144 29578
rect 29092 29514 29144 29520
rect 29000 26580 29052 26586
rect 29000 26522 29052 26528
rect 28906 25936 28962 25945
rect 28906 25871 28962 25880
rect 28920 24206 28948 25871
rect 29012 25294 29040 26522
rect 29000 25288 29052 25294
rect 29000 25230 29052 25236
rect 28908 24200 28960 24206
rect 28908 24142 28960 24148
rect 28356 23860 28408 23866
rect 28356 23802 28408 23808
rect 28264 23520 28316 23526
rect 28264 23462 28316 23468
rect 28276 23118 28304 23462
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 28356 22636 28408 22642
rect 28356 22578 28408 22584
rect 28368 22234 28396 22578
rect 28356 22228 28408 22234
rect 28356 22170 28408 22176
rect 28172 22160 28224 22166
rect 28172 22102 28224 22108
rect 29104 22094 29132 29514
rect 29288 29170 29316 29990
rect 29276 29164 29328 29170
rect 29276 29106 29328 29112
rect 29288 28626 29316 29106
rect 29276 28620 29328 28626
rect 29276 28562 29328 28568
rect 29288 28150 29316 28562
rect 29276 28144 29328 28150
rect 29276 28086 29328 28092
rect 29288 27538 29316 28086
rect 29380 27538 29408 31726
rect 29276 27532 29328 27538
rect 29276 27474 29328 27480
rect 29368 27532 29420 27538
rect 29368 27474 29420 27480
rect 29288 26994 29316 27474
rect 29276 26988 29328 26994
rect 29276 26930 29328 26936
rect 29288 26042 29316 26930
rect 29276 26036 29328 26042
rect 29276 25978 29328 25984
rect 29288 25362 29316 25978
rect 29276 25356 29328 25362
rect 29276 25298 29328 25304
rect 29288 24818 29316 25298
rect 29276 24812 29328 24818
rect 29276 24754 29328 24760
rect 29184 24744 29236 24750
rect 29184 24686 29236 24692
rect 29196 24410 29224 24686
rect 29184 24404 29236 24410
rect 29184 24346 29236 24352
rect 29276 23316 29328 23322
rect 29276 23258 29328 23264
rect 29104 22066 29224 22094
rect 28632 22024 28684 22030
rect 28632 21966 28684 21972
rect 28080 21888 28132 21894
rect 28080 21830 28132 21836
rect 28644 21690 28672 21966
rect 28632 21684 28684 21690
rect 28632 21626 28684 21632
rect 27252 21140 27304 21146
rect 27252 21082 27304 21088
rect 27988 21140 28040 21146
rect 27988 21082 28040 21088
rect 28356 20868 28408 20874
rect 28356 20810 28408 20816
rect 28368 20602 28396 20810
rect 28816 20800 28868 20806
rect 28816 20742 28868 20748
rect 28356 20596 28408 20602
rect 28356 20538 28408 20544
rect 28828 20262 28856 20742
rect 28816 20256 28868 20262
rect 28816 20198 28868 20204
rect 27160 19304 27212 19310
rect 27160 19246 27212 19252
rect 27080 16546 27292 16574
rect 26424 15632 26476 15638
rect 26424 15574 26476 15580
rect 26608 15496 26660 15502
rect 26528 15456 26608 15484
rect 26528 15366 26556 15456
rect 26608 15438 26660 15444
rect 26516 15360 26568 15366
rect 26516 15302 26568 15308
rect 26422 14648 26478 14657
rect 26422 14583 26424 14592
rect 26476 14583 26478 14592
rect 26424 14554 26476 14560
rect 26436 14346 26464 14554
rect 26608 14408 26660 14414
rect 26608 14350 26660 14356
rect 26424 14340 26476 14346
rect 26424 14282 26476 14288
rect 26344 12406 26464 12434
rect 26332 11824 26384 11830
rect 26332 11766 26384 11772
rect 26240 11076 26292 11082
rect 26240 11018 26292 11024
rect 26252 10577 26280 11018
rect 26238 10568 26294 10577
rect 26238 10503 26294 10512
rect 26344 8906 26372 11766
rect 26436 10470 26464 12406
rect 26620 12238 26648 14350
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 26424 10464 26476 10470
rect 26424 10406 26476 10412
rect 26436 9330 26464 10406
rect 26436 9302 26556 9330
rect 26422 9208 26478 9217
rect 26422 9143 26424 9152
rect 26476 9143 26478 9152
rect 26424 9114 26476 9120
rect 26332 8900 26384 8906
rect 26332 8842 26384 8848
rect 26238 8528 26294 8537
rect 26238 8463 26240 8472
rect 26292 8463 26294 8472
rect 26240 8434 26292 8440
rect 26148 8356 26200 8362
rect 26148 8298 26200 8304
rect 26240 7744 26292 7750
rect 26240 7686 26292 7692
rect 26252 7546 26280 7686
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 26146 6080 26202 6089
rect 26146 6015 26202 6024
rect 26160 5914 26188 6015
rect 26148 5908 26200 5914
rect 26148 5850 26200 5856
rect 25044 5636 25096 5642
rect 25044 5578 25096 5584
rect 24952 5296 25004 5302
rect 24952 5238 25004 5244
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 24584 4820 24636 4826
rect 24584 4762 24636 4768
rect 23848 4548 23900 4554
rect 23848 4490 23900 4496
rect 23572 4276 23624 4282
rect 23572 4218 23624 4224
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22848 2774 22876 3334
rect 23032 3194 23060 3674
rect 23216 3194 23244 3878
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 23492 3126 23520 4082
rect 23860 3534 23888 4490
rect 23940 4208 23992 4214
rect 24596 4185 24624 4762
rect 23940 4150 23992 4156
rect 24582 4176 24638 4185
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 23952 3466 23980 4150
rect 24216 4140 24268 4146
rect 24582 4111 24638 4120
rect 24216 4082 24268 4088
rect 24032 4072 24084 4078
rect 24032 4014 24084 4020
rect 23940 3460 23992 3466
rect 23940 3402 23992 3408
rect 23848 3392 23900 3398
rect 23848 3334 23900 3340
rect 23480 3120 23532 3126
rect 23480 3062 23532 3068
rect 22756 2746 22876 2774
rect 22468 2440 22520 2446
rect 22468 2382 22520 2388
rect 22756 800 22784 2746
rect 23296 2304 23348 2310
rect 23296 2246 23348 2252
rect 23308 800 23336 2246
rect 23860 800 23888 3334
rect 24044 3194 24072 4014
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 24124 3120 24176 3126
rect 24124 3062 24176 3068
rect 24136 2514 24164 3062
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 24228 2009 24256 4082
rect 24584 3528 24636 3534
rect 24768 3528 24820 3534
rect 24636 3476 24768 3482
rect 24584 3470 24820 3476
rect 24596 3454 24808 3470
rect 24952 3392 25004 3398
rect 24952 3334 25004 3340
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24596 2825 24624 2994
rect 24582 2816 24638 2825
rect 24582 2751 24638 2760
rect 24400 2576 24452 2582
rect 24400 2518 24452 2524
rect 24214 2000 24270 2009
rect 24214 1935 24270 1944
rect 24412 800 24440 2518
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 24504 2106 24532 2246
rect 24492 2100 24544 2106
rect 24492 2042 24544 2048
rect 24964 800 24992 3334
rect 25056 2446 25084 5578
rect 26528 5302 26556 9302
rect 25596 5296 25648 5302
rect 25596 5238 25648 5244
rect 26332 5296 26384 5302
rect 26332 5238 26384 5244
rect 26516 5296 26568 5302
rect 26516 5238 26568 5244
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 25516 3505 25544 3878
rect 25608 3534 25636 5238
rect 26240 4004 26292 4010
rect 26240 3946 26292 3952
rect 25870 3632 25926 3641
rect 26252 3602 26280 3946
rect 25870 3567 25926 3576
rect 26240 3596 26292 3602
rect 25596 3528 25648 3534
rect 25502 3496 25558 3505
rect 25596 3470 25648 3476
rect 25502 3431 25558 3440
rect 25884 3194 25912 3567
rect 26240 3538 26292 3544
rect 25872 3188 25924 3194
rect 25872 3130 25924 3136
rect 25504 2508 25556 2514
rect 25504 2450 25556 2456
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 25516 800 25544 2450
rect 26344 2446 26372 5238
rect 26422 5128 26478 5137
rect 26422 5063 26478 5072
rect 26436 4554 26464 5063
rect 26424 4548 26476 4554
rect 26424 4490 26476 4496
rect 26424 3732 26476 3738
rect 26424 3674 26476 3680
rect 26436 3602 26464 3674
rect 26896 3602 26924 16546
rect 27160 13320 27212 13326
rect 27160 13262 27212 13268
rect 27172 12918 27200 13262
rect 27160 12912 27212 12918
rect 27160 12854 27212 12860
rect 27172 12306 27200 12854
rect 27264 12714 27292 16546
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27436 14000 27488 14006
rect 27436 13942 27488 13948
rect 27252 12708 27304 12714
rect 27252 12650 27304 12656
rect 27160 12300 27212 12306
rect 27160 12242 27212 12248
rect 27172 11830 27200 12242
rect 27160 11824 27212 11830
rect 27160 11766 27212 11772
rect 27172 11218 27200 11766
rect 27160 11212 27212 11218
rect 27160 11154 27212 11160
rect 27172 10674 27200 11154
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 27172 10266 27200 10610
rect 27160 10260 27212 10266
rect 27160 10202 27212 10208
rect 26976 9376 27028 9382
rect 26976 9318 27028 9324
rect 26988 8838 27016 9318
rect 26976 8832 27028 8838
rect 26976 8774 27028 8780
rect 27264 4706 27292 12650
rect 27448 12434 27476 13942
rect 27356 12406 27476 12434
rect 27356 9178 27384 12406
rect 27540 10996 27568 15302
rect 28540 14816 28592 14822
rect 28540 14758 28592 14764
rect 28552 14414 28580 14758
rect 28540 14408 28592 14414
rect 28540 14350 28592 14356
rect 27710 12200 27766 12209
rect 27710 12135 27712 12144
rect 27764 12135 27766 12144
rect 27712 12106 27764 12112
rect 27620 11756 27672 11762
rect 27620 11698 27672 11704
rect 27448 10968 27568 10996
rect 27448 9382 27476 10968
rect 27632 10606 27660 11698
rect 28356 10668 28408 10674
rect 28356 10610 28408 10616
rect 27620 10600 27672 10606
rect 27620 10542 27672 10548
rect 28368 9586 28396 10610
rect 28356 9580 28408 9586
rect 28356 9522 28408 9528
rect 27436 9376 27488 9382
rect 27436 9318 27488 9324
rect 27344 9172 27396 9178
rect 27344 9114 27396 9120
rect 27356 5642 27384 9114
rect 28368 8906 28396 9522
rect 28356 8900 28408 8906
rect 28356 8842 28408 8848
rect 28368 8498 28396 8842
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 27436 8288 27488 8294
rect 27436 8230 27488 8236
rect 27344 5636 27396 5642
rect 27344 5578 27396 5584
rect 26988 4678 27292 4706
rect 26988 4010 27016 4678
rect 27068 4616 27120 4622
rect 27068 4558 27120 4564
rect 27080 4078 27108 4558
rect 27160 4480 27212 4486
rect 27160 4422 27212 4428
rect 27172 4146 27200 4422
rect 27160 4140 27212 4146
rect 27160 4082 27212 4088
rect 27068 4072 27120 4078
rect 27068 4014 27120 4020
rect 26976 4004 27028 4010
rect 26976 3946 27028 3952
rect 27080 3738 27108 4014
rect 27068 3732 27120 3738
rect 27068 3674 27120 3680
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 26884 3596 26936 3602
rect 26884 3538 26936 3544
rect 27160 3596 27212 3602
rect 27160 3538 27212 3544
rect 26896 2922 26924 3538
rect 26884 2916 26936 2922
rect 26884 2858 26936 2864
rect 26516 2644 26568 2650
rect 26516 2586 26568 2592
rect 26608 2644 26660 2650
rect 26608 2586 26660 2592
rect 26332 2440 26384 2446
rect 26332 2382 26384 2388
rect 26056 2304 26108 2310
rect 26056 2246 26108 2252
rect 26068 800 26096 2246
rect 26528 2106 26556 2586
rect 26516 2100 26568 2106
rect 26516 2042 26568 2048
rect 26620 800 26648 2586
rect 27172 800 27200 3538
rect 27448 3126 27476 8230
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 27632 6798 27660 7822
rect 27620 6792 27672 6798
rect 27620 6734 27672 6740
rect 28356 6792 28408 6798
rect 28356 6734 28408 6740
rect 28368 6390 28396 6734
rect 28828 6458 28856 20198
rect 29196 20058 29224 22066
rect 29184 20052 29236 20058
rect 29184 19994 29236 20000
rect 29184 19168 29236 19174
rect 29184 19110 29236 19116
rect 29196 11898 29224 19110
rect 29288 12434 29316 23258
rect 29368 21344 29420 21350
rect 29368 21286 29420 21292
rect 29380 21078 29408 21286
rect 29368 21072 29420 21078
rect 29368 21014 29420 21020
rect 29472 20942 29500 36178
rect 30012 36168 30064 36174
rect 30012 36110 30064 36116
rect 30024 35630 30052 36110
rect 30012 35624 30064 35630
rect 30012 35566 30064 35572
rect 30024 35086 30052 35566
rect 30116 35494 30144 37130
rect 30196 36712 30248 36718
rect 30196 36654 30248 36660
rect 30208 36174 30236 36654
rect 30196 36168 30248 36174
rect 30196 36110 30248 36116
rect 30286 36136 30342 36145
rect 30286 36071 30288 36080
rect 30340 36071 30342 36080
rect 30288 36042 30340 36048
rect 30392 35834 30420 37198
rect 30484 36922 30512 39200
rect 31036 39114 31064 39200
rect 31128 39114 31156 39222
rect 31036 39086 31156 39114
rect 31116 37256 31168 37262
rect 31116 37198 31168 37204
rect 30472 36916 30524 36922
rect 30472 36858 30524 36864
rect 30380 35828 30432 35834
rect 30380 35770 30432 35776
rect 31128 35494 31156 37198
rect 31404 37126 31432 39222
rect 31574 39200 31630 40000
rect 32126 39200 32182 40000
rect 32232 39222 32536 39250
rect 31588 37194 31616 39200
rect 32140 39114 32168 39200
rect 32232 39114 32260 39222
rect 32140 39086 32260 39114
rect 32508 37262 32536 39222
rect 32678 39200 32734 40000
rect 33230 39200 33286 40000
rect 33782 39200 33838 40000
rect 34334 39200 34390 40000
rect 34886 39200 34942 40000
rect 34992 39222 35388 39250
rect 32220 37256 32272 37262
rect 32220 37198 32272 37204
rect 32404 37256 32456 37262
rect 32404 37198 32456 37204
rect 32496 37256 32548 37262
rect 32496 37198 32548 37204
rect 31576 37188 31628 37194
rect 31576 37130 31628 37136
rect 31392 37120 31444 37126
rect 31392 37062 31444 37068
rect 31300 36780 31352 36786
rect 31300 36722 31352 36728
rect 30104 35488 30156 35494
rect 30104 35430 30156 35436
rect 31116 35488 31168 35494
rect 31116 35430 31168 35436
rect 30012 35080 30064 35086
rect 30012 35022 30064 35028
rect 30024 34678 30052 35022
rect 29644 34672 29696 34678
rect 29644 34614 29696 34620
rect 30012 34672 30064 34678
rect 30012 34614 30064 34620
rect 29656 34066 29684 34614
rect 29644 34060 29696 34066
rect 29644 34002 29696 34008
rect 29656 33318 29684 34002
rect 29644 33312 29696 33318
rect 29644 33254 29696 33260
rect 29656 32366 29684 33254
rect 29736 32428 29788 32434
rect 29736 32370 29788 32376
rect 29644 32360 29696 32366
rect 29644 32302 29696 32308
rect 29552 32020 29604 32026
rect 29552 31962 29604 31968
rect 29564 29617 29592 31962
rect 29656 31414 29684 32302
rect 29748 32026 29776 32370
rect 29736 32020 29788 32026
rect 29736 31962 29788 31968
rect 29644 31408 29696 31414
rect 29644 31350 29696 31356
rect 29550 29608 29606 29617
rect 29550 29543 29606 29552
rect 29736 28076 29788 28082
rect 29736 28018 29788 28024
rect 29552 24812 29604 24818
rect 29552 24754 29604 24760
rect 29564 24410 29592 24754
rect 29748 24682 29776 28018
rect 30116 27606 30144 35430
rect 30196 34604 30248 34610
rect 30196 34546 30248 34552
rect 30208 34202 30236 34546
rect 30196 34196 30248 34202
rect 30196 34138 30248 34144
rect 31022 32328 31078 32337
rect 31022 32263 31024 32272
rect 31076 32263 31078 32272
rect 31024 32234 31076 32240
rect 30656 31680 30708 31686
rect 30656 31622 30708 31628
rect 30288 30048 30340 30054
rect 30288 29990 30340 29996
rect 30300 29850 30328 29990
rect 30288 29844 30340 29850
rect 30288 29786 30340 29792
rect 30564 29164 30616 29170
rect 30564 29106 30616 29112
rect 30104 27600 30156 27606
rect 30104 27542 30156 27548
rect 29736 24676 29788 24682
rect 29736 24618 29788 24624
rect 29828 24608 29880 24614
rect 29828 24550 29880 24556
rect 29552 24404 29604 24410
rect 29552 24346 29604 24352
rect 29840 24206 29868 24550
rect 29828 24200 29880 24206
rect 29656 24148 29828 24154
rect 29656 24142 29880 24148
rect 30012 24200 30064 24206
rect 30012 24142 30064 24148
rect 29656 24126 29868 24142
rect 29552 23724 29604 23730
rect 29552 23666 29604 23672
rect 29564 23322 29592 23666
rect 29656 23662 29684 24126
rect 29644 23656 29696 23662
rect 29644 23598 29696 23604
rect 29552 23316 29604 23322
rect 29552 23258 29604 23264
rect 29656 23186 29684 23598
rect 29644 23180 29696 23186
rect 29644 23122 29696 23128
rect 30024 22778 30052 24142
rect 30012 22772 30064 22778
rect 30012 22714 30064 22720
rect 29828 22636 29880 22642
rect 29828 22578 29880 22584
rect 29644 21344 29696 21350
rect 29644 21286 29696 21292
rect 29460 20936 29512 20942
rect 29460 20878 29512 20884
rect 29550 13288 29606 13297
rect 29550 13223 29606 13232
rect 29564 12918 29592 13223
rect 29552 12912 29604 12918
rect 29552 12854 29604 12860
rect 29288 12406 29500 12434
rect 29184 11892 29236 11898
rect 29184 11834 29236 11840
rect 29276 9376 29328 9382
rect 29368 9376 29420 9382
rect 29276 9318 29328 9324
rect 29366 9344 29368 9353
rect 29420 9344 29422 9353
rect 29184 9172 29236 9178
rect 29184 9114 29236 9120
rect 29092 7812 29144 7818
rect 29092 7754 29144 7760
rect 29104 7546 29132 7754
rect 29092 7540 29144 7546
rect 29092 7482 29144 7488
rect 28816 6452 28868 6458
rect 28816 6394 28868 6400
rect 28356 6384 28408 6390
rect 28356 6326 28408 6332
rect 28998 6352 29054 6361
rect 27618 5808 27674 5817
rect 27618 5743 27674 5752
rect 27632 5710 27660 5743
rect 28368 5710 28396 6326
rect 28998 6287 29000 6296
rect 29052 6287 29054 6296
rect 29000 6258 29052 6264
rect 29196 5846 29224 9114
rect 29288 8634 29316 9318
rect 29366 9279 29422 9288
rect 29276 8628 29328 8634
rect 29276 8570 29328 8576
rect 29184 5840 29236 5846
rect 29184 5782 29236 5788
rect 27620 5704 27672 5710
rect 27620 5646 27672 5652
rect 28356 5704 28408 5710
rect 28356 5646 28408 5652
rect 27712 5296 27764 5302
rect 27712 5238 27764 5244
rect 27436 3120 27488 3126
rect 27436 3062 27488 3068
rect 27724 1873 27752 5238
rect 27804 5228 27856 5234
rect 27804 5170 27856 5176
rect 27816 3534 27844 5170
rect 28368 5166 28396 5646
rect 29196 5642 29224 5782
rect 29184 5636 29236 5642
rect 29184 5578 29236 5584
rect 28356 5160 28408 5166
rect 28356 5102 28408 5108
rect 28368 4622 28396 5102
rect 28724 5024 28776 5030
rect 28724 4966 28776 4972
rect 29368 5024 29420 5030
rect 29368 4966 29420 4972
rect 28356 4616 28408 4622
rect 28356 4558 28408 4564
rect 28264 4140 28316 4146
rect 28264 4082 28316 4088
rect 28078 3768 28134 3777
rect 28078 3703 28134 3712
rect 27804 3528 27856 3534
rect 27804 3470 27856 3476
rect 28092 3126 28120 3703
rect 28080 3120 28132 3126
rect 28080 3062 28132 3068
rect 28080 2372 28132 2378
rect 28080 2314 28132 2320
rect 27710 1864 27766 1873
rect 27710 1799 27766 1808
rect 27724 870 27844 898
rect 27724 800 27752 870
rect 1766 0 1822 800
rect 2318 0 2374 800
rect 2870 0 2926 800
rect 3422 0 3478 800
rect 3974 0 4030 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5630 0 5686 800
rect 6182 0 6238 800
rect 6734 0 6790 800
rect 7286 0 7342 800
rect 7838 0 7894 800
rect 8390 0 8446 800
rect 8942 0 8998 800
rect 9494 0 9550 800
rect 10046 0 10102 800
rect 10598 0 10654 800
rect 11150 0 11206 800
rect 11702 0 11758 800
rect 12254 0 12310 800
rect 12806 0 12862 800
rect 13358 0 13414 800
rect 13910 0 13966 800
rect 14462 0 14518 800
rect 15014 0 15070 800
rect 15566 0 15622 800
rect 16118 0 16174 800
rect 16670 0 16726 800
rect 17222 0 17278 800
rect 17774 0 17830 800
rect 18326 0 18382 800
rect 18878 0 18934 800
rect 19430 0 19486 800
rect 19982 0 20038 800
rect 20534 0 20590 800
rect 21086 0 21142 800
rect 21638 0 21694 800
rect 22190 0 22246 800
rect 22742 0 22798 800
rect 23294 0 23350 800
rect 23846 0 23902 800
rect 24398 0 24454 800
rect 24950 0 25006 800
rect 25502 0 25558 800
rect 26054 0 26110 800
rect 26606 0 26662 800
rect 27158 0 27214 800
rect 27710 0 27766 800
rect 27816 762 27844 870
rect 28092 762 28120 2314
rect 28276 800 28304 4082
rect 28368 4060 28396 4558
rect 28446 4312 28502 4321
rect 28502 4256 28580 4264
rect 28446 4247 28448 4256
rect 28500 4236 28580 4256
rect 28448 4218 28500 4224
rect 28448 4072 28500 4078
rect 28368 4032 28448 4060
rect 28368 3058 28396 4032
rect 28448 4014 28500 4020
rect 28552 3942 28580 4236
rect 28540 3936 28592 3942
rect 28540 3878 28592 3884
rect 28448 3664 28500 3670
rect 28448 3606 28500 3612
rect 28460 3398 28488 3606
rect 28448 3392 28500 3398
rect 28448 3334 28500 3340
rect 28356 3052 28408 3058
rect 28356 2994 28408 3000
rect 28736 2446 28764 4966
rect 29000 4480 29052 4486
rect 29000 4422 29052 4428
rect 29012 4146 29040 4422
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 28998 3768 29054 3777
rect 28998 3703 29000 3712
rect 29052 3703 29054 3712
rect 29092 3732 29144 3738
rect 29000 3674 29052 3680
rect 29092 3674 29144 3680
rect 29012 2582 29040 3674
rect 29000 2576 29052 2582
rect 29000 2518 29052 2524
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 28828 2378 29040 2394
rect 28828 2372 29052 2378
rect 28828 2366 29000 2372
rect 28828 800 28856 2366
rect 29000 2314 29052 2320
rect 29104 2310 29132 3674
rect 29380 2446 29408 4966
rect 29472 3942 29500 12406
rect 29656 5710 29684 21286
rect 29840 20602 29868 22578
rect 30012 22024 30064 22030
rect 30012 21966 30064 21972
rect 30024 21146 30052 21966
rect 30116 21962 30144 27542
rect 30196 27532 30248 27538
rect 30196 27474 30248 27480
rect 30208 23798 30236 27474
rect 30472 27328 30524 27334
rect 30472 27270 30524 27276
rect 30380 26376 30432 26382
rect 30380 26318 30432 26324
rect 30392 25974 30420 26318
rect 30380 25968 30432 25974
rect 30380 25910 30432 25916
rect 30196 23792 30248 23798
rect 30196 23734 30248 23740
rect 30208 23322 30236 23734
rect 30196 23316 30248 23322
rect 30196 23258 30248 23264
rect 30380 23112 30432 23118
rect 30380 23054 30432 23060
rect 30196 22636 30248 22642
rect 30196 22578 30248 22584
rect 30208 22098 30236 22578
rect 30392 22574 30420 23054
rect 30380 22568 30432 22574
rect 30380 22510 30432 22516
rect 30392 22166 30420 22510
rect 30484 22506 30512 27270
rect 30576 22710 30604 29106
rect 30668 27470 30696 31622
rect 30656 27464 30708 27470
rect 30656 27406 30708 27412
rect 30748 27396 30800 27402
rect 30748 27338 30800 27344
rect 30656 26784 30708 26790
rect 30656 26726 30708 26732
rect 30668 25158 30696 26726
rect 30656 25152 30708 25158
rect 30656 25094 30708 25100
rect 30656 23724 30708 23730
rect 30656 23666 30708 23672
rect 30564 22704 30616 22710
rect 30564 22646 30616 22652
rect 30472 22500 30524 22506
rect 30472 22442 30524 22448
rect 30380 22160 30432 22166
rect 30380 22102 30432 22108
rect 30196 22092 30248 22098
rect 30196 22034 30248 22040
rect 30288 22092 30340 22098
rect 30288 22034 30340 22040
rect 30300 21978 30328 22034
rect 30104 21956 30156 21962
rect 30104 21898 30156 21904
rect 30208 21950 30328 21978
rect 30208 21486 30236 21950
rect 30196 21480 30248 21486
rect 30196 21422 30248 21428
rect 30012 21140 30064 21146
rect 30012 21082 30064 21088
rect 30208 21010 30236 21422
rect 30196 21004 30248 21010
rect 30196 20946 30248 20952
rect 30104 20936 30156 20942
rect 30104 20878 30156 20884
rect 30116 20602 30144 20878
rect 29828 20596 29880 20602
rect 29828 20538 29880 20544
rect 30104 20596 30156 20602
rect 30104 20538 30156 20544
rect 29920 20460 29972 20466
rect 29920 20402 29972 20408
rect 29932 20058 29960 20402
rect 30208 20398 30236 20946
rect 30012 20392 30064 20398
rect 30012 20334 30064 20340
rect 30196 20392 30248 20398
rect 30196 20334 30248 20340
rect 29920 20052 29972 20058
rect 29920 19994 29972 20000
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 29932 19174 29960 19790
rect 29920 19168 29972 19174
rect 29920 19110 29972 19116
rect 29736 17060 29788 17066
rect 29736 17002 29788 17008
rect 29748 12102 29776 17002
rect 29932 14890 29960 19110
rect 29920 14884 29972 14890
rect 29920 14826 29972 14832
rect 29736 12096 29788 12102
rect 29736 12038 29788 12044
rect 29644 5704 29696 5710
rect 29644 5646 29696 5652
rect 29748 5098 29776 12038
rect 30024 11218 30052 20334
rect 30564 19780 30616 19786
rect 30564 19722 30616 19728
rect 30104 19712 30156 19718
rect 30104 19654 30156 19660
rect 30116 19378 30144 19654
rect 30104 19372 30156 19378
rect 30104 19314 30156 19320
rect 30288 15632 30340 15638
rect 30288 15574 30340 15580
rect 30300 15026 30328 15574
rect 30288 15020 30340 15026
rect 30288 14962 30340 14968
rect 30196 14884 30248 14890
rect 30196 14826 30248 14832
rect 30104 13932 30156 13938
rect 30104 13874 30156 13880
rect 30116 13190 30144 13874
rect 30104 13184 30156 13190
rect 30104 13126 30156 13132
rect 30012 11212 30064 11218
rect 30012 11154 30064 11160
rect 29736 5092 29788 5098
rect 29736 5034 29788 5040
rect 29828 5024 29880 5030
rect 29828 4966 29880 4972
rect 29460 3936 29512 3942
rect 29460 3878 29512 3884
rect 29644 3120 29696 3126
rect 29644 3062 29696 3068
rect 29460 2848 29512 2854
rect 29460 2790 29512 2796
rect 29368 2440 29420 2446
rect 29368 2382 29420 2388
rect 29092 2304 29144 2310
rect 29472 2292 29500 2790
rect 29092 2246 29144 2252
rect 29380 2264 29500 2292
rect 29552 2304 29604 2310
rect 29380 800 29408 2264
rect 29552 2246 29604 2252
rect 29564 1970 29592 2246
rect 29656 2106 29684 3062
rect 29840 2378 29868 4966
rect 29920 4480 29972 4486
rect 29920 4422 29972 4428
rect 29932 4214 29960 4422
rect 29920 4208 29972 4214
rect 29920 4150 29972 4156
rect 30116 3738 30144 13126
rect 30208 10810 30236 14826
rect 30472 14816 30524 14822
rect 30472 14758 30524 14764
rect 30288 14272 30340 14278
rect 30288 14214 30340 14220
rect 30300 13258 30328 14214
rect 30380 13796 30432 13802
rect 30380 13738 30432 13744
rect 30288 13252 30340 13258
rect 30288 13194 30340 13200
rect 30392 11354 30420 13738
rect 30484 12238 30512 14758
rect 30472 12232 30524 12238
rect 30472 12174 30524 12180
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 30196 10804 30248 10810
rect 30196 10746 30248 10752
rect 30472 10056 30524 10062
rect 30472 9998 30524 10004
rect 30484 8090 30512 9998
rect 30576 9874 30604 19722
rect 30668 19446 30696 23666
rect 30760 22506 30788 27338
rect 31128 27062 31156 35430
rect 31312 34950 31340 36722
rect 31852 36100 31904 36106
rect 31852 36042 31904 36048
rect 31668 36032 31720 36038
rect 31668 35974 31720 35980
rect 31392 35216 31444 35222
rect 31390 35184 31392 35193
rect 31444 35184 31446 35193
rect 31390 35119 31446 35128
rect 31300 34944 31352 34950
rect 31300 34886 31352 34892
rect 31208 31952 31260 31958
rect 31208 31894 31260 31900
rect 31116 27056 31168 27062
rect 31116 26998 31168 27004
rect 31220 26081 31248 31894
rect 31206 26072 31262 26081
rect 31206 26007 31262 26016
rect 30932 25152 30984 25158
rect 30932 25094 30984 25100
rect 31024 25152 31076 25158
rect 31024 25094 31076 25100
rect 30840 24132 30892 24138
rect 30840 24074 30892 24080
rect 30852 23730 30880 24074
rect 30944 23769 30972 25094
rect 31036 24954 31064 25094
rect 31024 24948 31076 24954
rect 31024 24890 31076 24896
rect 31208 24812 31260 24818
rect 31208 24754 31260 24760
rect 31024 24200 31076 24206
rect 31024 24142 31076 24148
rect 31036 23866 31064 24142
rect 31220 23866 31248 24754
rect 31024 23860 31076 23866
rect 31024 23802 31076 23808
rect 31208 23860 31260 23866
rect 31208 23802 31260 23808
rect 30930 23760 30986 23769
rect 30840 23724 30892 23730
rect 30930 23695 30986 23704
rect 31024 23724 31076 23730
rect 30840 23666 30892 23672
rect 31024 23666 31076 23672
rect 30852 22778 30880 23666
rect 30932 23112 30984 23118
rect 30932 23054 30984 23060
rect 30840 22772 30892 22778
rect 30840 22714 30892 22720
rect 30748 22500 30800 22506
rect 30748 22442 30800 22448
rect 30944 21146 30972 23054
rect 31036 21690 31064 23666
rect 31024 21684 31076 21690
rect 31024 21626 31076 21632
rect 30932 21140 30984 21146
rect 30932 21082 30984 21088
rect 31312 20942 31340 34886
rect 31680 34105 31708 35974
rect 31864 34785 31892 36042
rect 32232 35894 32260 37198
rect 32416 36174 32444 37198
rect 32404 36168 32456 36174
rect 32404 36110 32456 36116
rect 32140 35866 32260 35894
rect 32140 35494 32168 35866
rect 32692 35834 32720 39200
rect 33244 35834 33272 39200
rect 33796 37618 33824 39200
rect 33796 37590 33916 37618
rect 33784 36712 33836 36718
rect 33784 36654 33836 36660
rect 33796 36242 33824 36654
rect 33784 36236 33836 36242
rect 33784 36178 33836 36184
rect 32680 35828 32732 35834
rect 32680 35770 32732 35776
rect 33232 35828 33284 35834
rect 33232 35770 33284 35776
rect 32864 35556 32916 35562
rect 32864 35498 32916 35504
rect 32128 35488 32180 35494
rect 32128 35430 32180 35436
rect 31944 35012 31996 35018
rect 31944 34954 31996 34960
rect 31850 34776 31906 34785
rect 31850 34711 31906 34720
rect 31666 34096 31722 34105
rect 31666 34031 31722 34040
rect 31392 32020 31444 32026
rect 31392 31962 31444 31968
rect 31404 24682 31432 31962
rect 31852 29504 31904 29510
rect 31852 29446 31904 29452
rect 31760 28484 31812 28490
rect 31760 28426 31812 28432
rect 31772 27577 31800 28426
rect 31758 27568 31814 27577
rect 31758 27503 31814 27512
rect 31760 27464 31812 27470
rect 31760 27406 31812 27412
rect 31484 27124 31536 27130
rect 31484 27066 31536 27072
rect 31496 26382 31524 27066
rect 31668 27056 31720 27062
rect 31668 26998 31720 27004
rect 31484 26376 31536 26382
rect 31484 26318 31536 26324
rect 31392 24676 31444 24682
rect 31392 24618 31444 24624
rect 31576 24608 31628 24614
rect 31576 24550 31628 24556
rect 31588 24206 31616 24550
rect 31576 24200 31628 24206
rect 31576 24142 31628 24148
rect 31484 22160 31536 22166
rect 31484 22102 31536 22108
rect 31392 21616 31444 21622
rect 31392 21558 31444 21564
rect 31300 20936 31352 20942
rect 31300 20878 31352 20884
rect 30748 20800 30800 20806
rect 30748 20742 30800 20748
rect 30760 20262 30788 20742
rect 30748 20256 30800 20262
rect 30748 20198 30800 20204
rect 30656 19440 30708 19446
rect 30656 19382 30708 19388
rect 30760 16574 30788 20198
rect 31404 16574 31432 21558
rect 31496 21486 31524 22102
rect 31484 21480 31536 21486
rect 31484 21422 31536 21428
rect 31680 20874 31708 26998
rect 31772 23322 31800 27406
rect 31760 23316 31812 23322
rect 31760 23258 31812 23264
rect 31864 23050 31892 29446
rect 31956 27470 31984 34954
rect 32140 30938 32168 35430
rect 32128 30932 32180 30938
rect 32128 30874 32180 30880
rect 32140 30682 32168 30874
rect 32312 30728 32364 30734
rect 32140 30654 32260 30682
rect 32312 30670 32364 30676
rect 32128 30592 32180 30598
rect 32128 30534 32180 30540
rect 32036 27872 32088 27878
rect 32036 27814 32088 27820
rect 31944 27464 31996 27470
rect 31944 27406 31996 27412
rect 31944 26444 31996 26450
rect 31944 26386 31996 26392
rect 31956 25158 31984 26386
rect 31944 25152 31996 25158
rect 31944 25094 31996 25100
rect 32048 24206 32076 27814
rect 32140 24970 32168 30534
rect 32232 25106 32260 30654
rect 32324 29714 32352 30670
rect 32312 29708 32364 29714
rect 32312 29650 32364 29656
rect 32324 29238 32352 29650
rect 32312 29232 32364 29238
rect 32312 29174 32364 29180
rect 32324 28626 32352 29174
rect 32876 29034 32904 35498
rect 33796 35086 33824 36178
rect 33888 35834 33916 37590
rect 34244 37324 34296 37330
rect 34244 37266 34296 37272
rect 33968 36576 34020 36582
rect 33968 36518 34020 36524
rect 33980 36417 34008 36518
rect 33966 36408 34022 36417
rect 33966 36343 34022 36352
rect 33876 35828 33928 35834
rect 33876 35770 33928 35776
rect 33508 35080 33560 35086
rect 33508 35022 33560 35028
rect 33784 35080 33836 35086
rect 33784 35022 33836 35028
rect 33520 34406 33548 35022
rect 33048 34400 33100 34406
rect 33048 34342 33100 34348
rect 33140 34400 33192 34406
rect 33140 34342 33192 34348
rect 33508 34400 33560 34406
rect 33508 34342 33560 34348
rect 33060 33561 33088 34342
rect 33152 33862 33180 34342
rect 33232 33924 33284 33930
rect 33232 33866 33284 33872
rect 33140 33856 33192 33862
rect 33140 33798 33192 33804
rect 33046 33552 33102 33561
rect 33046 33487 33102 33496
rect 33152 32910 33180 33798
rect 33244 33522 33272 33866
rect 33232 33516 33284 33522
rect 33232 33458 33284 33464
rect 33140 32904 33192 32910
rect 33140 32846 33192 32852
rect 33152 31822 33180 32846
rect 33140 31816 33192 31822
rect 33140 31758 33192 31764
rect 33152 31346 33180 31758
rect 33140 31340 33192 31346
rect 33140 31282 33192 31288
rect 33140 31136 33192 31142
rect 33244 31124 33272 33458
rect 33322 32872 33378 32881
rect 33322 32807 33324 32816
rect 33376 32807 33378 32816
rect 33324 32778 33376 32784
rect 33192 31096 33272 31124
rect 33140 31078 33192 31084
rect 32864 29028 32916 29034
rect 32864 28970 32916 28976
rect 32312 28620 32364 28626
rect 32312 28562 32364 28568
rect 32324 27470 32352 28562
rect 32312 27464 32364 27470
rect 32312 27406 32364 27412
rect 32312 26444 32364 26450
rect 32312 26386 32364 26392
rect 32324 25974 32352 26386
rect 32312 25968 32364 25974
rect 32312 25910 32364 25916
rect 32324 25226 32352 25910
rect 32312 25220 32364 25226
rect 32312 25162 32364 25168
rect 32232 25078 32352 25106
rect 32140 24942 32260 24970
rect 32128 24812 32180 24818
rect 32128 24754 32180 24760
rect 32140 24410 32168 24754
rect 32128 24404 32180 24410
rect 32128 24346 32180 24352
rect 32232 24342 32260 24942
rect 32220 24336 32272 24342
rect 32220 24278 32272 24284
rect 32036 24200 32088 24206
rect 32036 24142 32088 24148
rect 31852 23044 31904 23050
rect 31852 22986 31904 22992
rect 32324 22930 32352 25078
rect 32680 24064 32732 24070
rect 32680 24006 32732 24012
rect 32692 23730 32720 24006
rect 32680 23724 32732 23730
rect 32680 23666 32732 23672
rect 32496 23656 32548 23662
rect 32496 23598 32548 23604
rect 32508 23322 32536 23598
rect 32496 23316 32548 23322
rect 32496 23258 32548 23264
rect 32508 23118 32536 23258
rect 32496 23112 32548 23118
rect 32496 23054 32548 23060
rect 32232 22902 32352 22930
rect 31668 20868 31720 20874
rect 31668 20810 31720 20816
rect 32232 20058 32260 22902
rect 32310 22808 32366 22817
rect 32508 22778 32536 23054
rect 32310 22743 32312 22752
rect 32364 22743 32366 22752
rect 32496 22772 32548 22778
rect 32312 22714 32364 22720
rect 32496 22714 32548 22720
rect 32772 21888 32824 21894
rect 32772 21830 32824 21836
rect 32784 21350 32812 21830
rect 32876 21554 32904 28970
rect 33048 27464 33100 27470
rect 33048 27406 33100 27412
rect 33060 27062 33088 27406
rect 33048 27056 33100 27062
rect 33048 26998 33100 27004
rect 33060 26450 33088 26998
rect 33048 26444 33100 26450
rect 33048 26386 33100 26392
rect 33152 26314 33180 31078
rect 33416 30252 33468 30258
rect 33416 30194 33468 30200
rect 33232 26988 33284 26994
rect 33232 26930 33284 26936
rect 33244 26602 33272 26930
rect 33244 26574 33364 26602
rect 33232 26512 33284 26518
rect 33232 26454 33284 26460
rect 33140 26308 33192 26314
rect 33140 26250 33192 26256
rect 33140 24812 33192 24818
rect 33140 24754 33192 24760
rect 33152 23866 33180 24754
rect 33244 24682 33272 26454
rect 33232 24676 33284 24682
rect 33232 24618 33284 24624
rect 33336 24426 33364 26574
rect 33428 26518 33456 30194
rect 33508 30048 33560 30054
rect 33508 29990 33560 29996
rect 33520 29850 33548 29990
rect 33508 29844 33560 29850
rect 33508 29786 33560 29792
rect 33416 26512 33468 26518
rect 33416 26454 33468 26460
rect 33416 26376 33468 26382
rect 33416 26318 33468 26324
rect 33428 25906 33456 26318
rect 33416 25900 33468 25906
rect 33416 25842 33468 25848
rect 33692 25288 33744 25294
rect 33692 25230 33744 25236
rect 33600 24608 33652 24614
rect 33600 24550 33652 24556
rect 33244 24398 33364 24426
rect 33244 24274 33272 24398
rect 33232 24268 33284 24274
rect 33232 24210 33284 24216
rect 33612 24070 33640 24550
rect 33600 24064 33652 24070
rect 33600 24006 33652 24012
rect 33140 23860 33192 23866
rect 33140 23802 33192 23808
rect 33140 23112 33192 23118
rect 33140 23054 33192 23060
rect 33152 22234 33180 23054
rect 33140 22228 33192 22234
rect 33140 22170 33192 22176
rect 32864 21548 32916 21554
rect 32864 21490 32916 21496
rect 32772 21344 32824 21350
rect 32772 21286 32824 21292
rect 32312 20800 32364 20806
rect 32312 20742 32364 20748
rect 32220 20052 32272 20058
rect 32220 19994 32272 20000
rect 30760 16546 30880 16574
rect 30656 15700 30708 15706
rect 30656 15642 30708 15648
rect 30668 11082 30696 15642
rect 30748 11212 30800 11218
rect 30748 11154 30800 11160
rect 30656 11076 30708 11082
rect 30656 11018 30708 11024
rect 30576 9846 30696 9874
rect 30564 9716 30616 9722
rect 30564 9658 30616 9664
rect 30576 8974 30604 9658
rect 30668 9178 30696 9846
rect 30656 9172 30708 9178
rect 30656 9114 30708 9120
rect 30564 8968 30616 8974
rect 30564 8910 30616 8916
rect 30668 8362 30696 9114
rect 30656 8356 30708 8362
rect 30656 8298 30708 8304
rect 30472 8084 30524 8090
rect 30472 8026 30524 8032
rect 30380 7472 30432 7478
rect 30378 7440 30380 7449
rect 30432 7440 30434 7449
rect 30288 7404 30340 7410
rect 30378 7375 30434 7384
rect 30288 7346 30340 7352
rect 30300 6458 30328 7346
rect 30760 6866 30788 11154
rect 30852 8090 30880 16546
rect 31220 16546 31432 16574
rect 32324 16574 32352 20742
rect 32680 19508 32732 19514
rect 32680 19450 32732 19456
rect 32324 16546 32536 16574
rect 30840 8084 30892 8090
rect 30840 8026 30892 8032
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30748 6860 30800 6866
rect 30748 6802 30800 6808
rect 30288 6452 30340 6458
rect 30288 6394 30340 6400
rect 30576 6390 30604 6802
rect 30840 6656 30892 6662
rect 30840 6598 30892 6604
rect 30564 6384 30616 6390
rect 30564 6326 30616 6332
rect 30656 6316 30708 6322
rect 30656 6258 30708 6264
rect 30564 5024 30616 5030
rect 30564 4966 30616 4972
rect 30104 3732 30156 3738
rect 30104 3674 30156 3680
rect 30196 3392 30248 3398
rect 30196 3334 30248 3340
rect 30208 3126 30236 3334
rect 30196 3120 30248 3126
rect 30196 3062 30248 3068
rect 30576 3058 30604 4966
rect 30104 3052 30156 3058
rect 30104 2994 30156 3000
rect 30564 3052 30616 3058
rect 30564 2994 30616 3000
rect 30116 2774 30144 2994
rect 30472 2848 30524 2854
rect 30472 2790 30524 2796
rect 29932 2746 30144 2774
rect 29828 2372 29880 2378
rect 29828 2314 29880 2320
rect 29644 2100 29696 2106
rect 29644 2042 29696 2048
rect 29552 1964 29604 1970
rect 29552 1906 29604 1912
rect 29932 800 29960 2746
rect 30484 800 30512 2790
rect 30668 2650 30696 6258
rect 30852 3194 30880 6598
rect 31220 4554 31248 16546
rect 32128 15496 32180 15502
rect 32128 15438 32180 15444
rect 32140 15026 32168 15438
rect 32128 15020 32180 15026
rect 32128 14962 32180 14968
rect 31852 14272 31904 14278
rect 31852 14214 31904 14220
rect 31864 14074 31892 14214
rect 31852 14068 31904 14074
rect 31852 14010 31904 14016
rect 31760 13320 31812 13326
rect 31760 13262 31812 13268
rect 31772 12782 31800 13262
rect 32140 12986 32168 14962
rect 32128 12980 32180 12986
rect 32128 12922 32180 12928
rect 31760 12776 31812 12782
rect 31760 12718 31812 12724
rect 31772 12238 31800 12718
rect 31760 12232 31812 12238
rect 31760 12174 31812 12180
rect 31944 12232 31996 12238
rect 31944 12174 31996 12180
rect 31760 11892 31812 11898
rect 31760 11834 31812 11840
rect 31484 7336 31536 7342
rect 31484 7278 31536 7284
rect 31300 7200 31352 7206
rect 31300 7142 31352 7148
rect 31208 4548 31260 4554
rect 31208 4490 31260 4496
rect 31220 4282 31248 4490
rect 31208 4276 31260 4282
rect 31208 4218 31260 4224
rect 30840 3188 30892 3194
rect 30840 3130 30892 3136
rect 31024 3052 31076 3058
rect 31024 2994 31076 3000
rect 30656 2644 30708 2650
rect 30656 2586 30708 2592
rect 31036 800 31064 2994
rect 31312 2922 31340 7142
rect 31496 6798 31524 7278
rect 31484 6792 31536 6798
rect 31484 6734 31536 6740
rect 31392 6452 31444 6458
rect 31392 6394 31444 6400
rect 31404 5914 31432 6394
rect 31392 5908 31444 5914
rect 31392 5850 31444 5856
rect 31496 5710 31524 6734
rect 31484 5704 31536 5710
rect 31484 5646 31536 5652
rect 31496 3398 31524 5646
rect 31576 5024 31628 5030
rect 31576 4966 31628 4972
rect 31588 4690 31616 4966
rect 31576 4684 31628 4690
rect 31576 4626 31628 4632
rect 31484 3392 31536 3398
rect 31484 3334 31536 3340
rect 31496 2990 31524 3334
rect 31484 2984 31536 2990
rect 31484 2926 31536 2932
rect 31300 2916 31352 2922
rect 31300 2858 31352 2864
rect 31312 2446 31340 2858
rect 31300 2440 31352 2446
rect 31300 2382 31352 2388
rect 31588 800 31616 4626
rect 31668 4276 31720 4282
rect 31668 4218 31720 4224
rect 31680 2650 31708 4218
rect 31772 3777 31800 11834
rect 31956 11150 31984 12174
rect 31944 11144 31996 11150
rect 31944 11086 31996 11092
rect 31956 9926 31984 11086
rect 31944 9920 31996 9926
rect 31944 9862 31996 9868
rect 31956 9586 31984 9862
rect 31944 9580 31996 9586
rect 31944 9522 31996 9528
rect 31956 8974 31984 9522
rect 31944 8968 31996 8974
rect 31944 8910 31996 8916
rect 32404 8968 32456 8974
rect 32404 8910 32456 8916
rect 32220 8288 32272 8294
rect 32220 8230 32272 8236
rect 32232 7886 32260 8230
rect 32416 7954 32444 8910
rect 32404 7948 32456 7954
rect 32404 7890 32456 7896
rect 32220 7880 32272 7886
rect 32220 7822 32272 7828
rect 32128 7404 32180 7410
rect 32128 7346 32180 7352
rect 32140 6662 32168 7346
rect 32312 7200 32364 7206
rect 32312 7142 32364 7148
rect 32324 6730 32352 7142
rect 32312 6724 32364 6730
rect 32312 6666 32364 6672
rect 32128 6656 32180 6662
rect 32128 6598 32180 6604
rect 32508 6458 32536 16546
rect 32588 14408 32640 14414
rect 32588 14350 32640 14356
rect 32600 11354 32628 14350
rect 32588 11348 32640 11354
rect 32588 11290 32640 11296
rect 32692 11082 32720 19450
rect 32784 16574 32812 21286
rect 33508 19304 33560 19310
rect 33508 19246 33560 19252
rect 33232 18080 33284 18086
rect 33232 18022 33284 18028
rect 32784 16546 32904 16574
rect 32680 11076 32732 11082
rect 32680 11018 32732 11024
rect 32772 7200 32824 7206
rect 32772 7142 32824 7148
rect 32496 6452 32548 6458
rect 32496 6394 32548 6400
rect 32036 6248 32088 6254
rect 32036 6190 32088 6196
rect 32048 5846 32076 6190
rect 32508 6118 32536 6394
rect 32496 6112 32548 6118
rect 32496 6054 32548 6060
rect 32036 5840 32088 5846
rect 32036 5782 32088 5788
rect 32048 4758 32076 5782
rect 32588 5636 32640 5642
rect 32588 5578 32640 5584
rect 32496 5568 32548 5574
rect 32496 5510 32548 5516
rect 32508 5166 32536 5510
rect 32496 5160 32548 5166
rect 32496 5102 32548 5108
rect 32036 4752 32088 4758
rect 32036 4694 32088 4700
rect 32048 4078 32076 4694
rect 32128 4616 32180 4622
rect 32128 4558 32180 4564
rect 32140 4282 32168 4558
rect 32128 4276 32180 4282
rect 32128 4218 32180 4224
rect 32496 4208 32548 4214
rect 32496 4150 32548 4156
rect 32036 4072 32088 4078
rect 32036 4014 32088 4020
rect 31758 3768 31814 3777
rect 31758 3703 31814 3712
rect 32220 3460 32272 3466
rect 32220 3402 32272 3408
rect 31760 3052 31812 3058
rect 31760 2994 31812 3000
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 31772 1737 31800 2994
rect 32128 2984 32180 2990
rect 32128 2926 32180 2932
rect 32140 2514 32168 2926
rect 32128 2508 32180 2514
rect 32128 2450 32180 2456
rect 31758 1728 31814 1737
rect 32232 1714 32260 3402
rect 32508 2582 32536 4150
rect 32600 4146 32628 5578
rect 32680 4616 32732 4622
rect 32680 4558 32732 4564
rect 32588 4140 32640 4146
rect 32588 4082 32640 4088
rect 32496 2576 32548 2582
rect 32496 2518 32548 2524
rect 31758 1663 31814 1672
rect 32140 1686 32260 1714
rect 32140 800 32168 1686
rect 32692 800 32720 4558
rect 32784 3126 32812 7142
rect 32876 5166 32904 16546
rect 33140 15496 33192 15502
rect 33140 15438 33192 15444
rect 33152 15162 33180 15438
rect 33140 15156 33192 15162
rect 33140 15098 33192 15104
rect 33244 9178 33272 18022
rect 33324 15428 33376 15434
rect 33324 15370 33376 15376
rect 33336 11286 33364 15370
rect 33416 14272 33468 14278
rect 33416 14214 33468 14220
rect 33428 12918 33456 14214
rect 33416 12912 33468 12918
rect 33416 12854 33468 12860
rect 33324 11280 33376 11286
rect 33324 11222 33376 11228
rect 33232 9172 33284 9178
rect 33232 9114 33284 9120
rect 33140 7744 33192 7750
rect 33140 7686 33192 7692
rect 32956 6180 33008 6186
rect 32956 6122 33008 6128
rect 32864 5160 32916 5166
rect 32864 5102 32916 5108
rect 32968 4622 32996 6122
rect 33152 5914 33180 7686
rect 33244 6390 33272 9114
rect 33416 7404 33468 7410
rect 33416 7346 33468 7352
rect 33232 6384 33284 6390
rect 33232 6326 33284 6332
rect 33244 5914 33272 6326
rect 33140 5908 33192 5914
rect 33140 5850 33192 5856
rect 33232 5908 33284 5914
rect 33232 5850 33284 5856
rect 33048 5092 33100 5098
rect 33048 5034 33100 5040
rect 33060 4690 33088 5034
rect 33048 4684 33100 4690
rect 33048 4626 33100 4632
rect 32956 4616 33008 4622
rect 32956 4558 33008 4564
rect 33060 4214 33088 4626
rect 33140 4480 33192 4486
rect 33140 4422 33192 4428
rect 33152 4282 33180 4422
rect 33140 4276 33192 4282
rect 33140 4218 33192 4224
rect 33048 4208 33100 4214
rect 33048 4150 33100 4156
rect 33232 4140 33284 4146
rect 33232 4082 33284 4088
rect 33048 4072 33100 4078
rect 33048 4014 33100 4020
rect 33060 3602 33088 4014
rect 33048 3596 33100 3602
rect 33048 3538 33100 3544
rect 32772 3120 32824 3126
rect 32772 3062 32824 3068
rect 33244 800 33272 4082
rect 33428 3398 33456 7346
rect 33416 3392 33468 3398
rect 33416 3334 33468 3340
rect 33520 3097 33548 19246
rect 33612 9110 33640 24006
rect 33704 22778 33732 25230
rect 33784 24676 33836 24682
rect 33784 24618 33836 24624
rect 33692 22772 33744 22778
rect 33692 22714 33744 22720
rect 33796 18426 33824 24618
rect 33784 18420 33836 18426
rect 33784 18362 33836 18368
rect 33692 14476 33744 14482
rect 33692 14418 33744 14424
rect 33704 11014 33732 14418
rect 33796 12986 33824 18362
rect 33980 17338 34008 36343
rect 34256 36174 34284 37266
rect 34348 36904 34376 39200
rect 34900 39114 34928 39200
rect 34992 39114 35020 39222
rect 34900 39086 35020 39114
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35072 37392 35124 37398
rect 35072 37334 35124 37340
rect 34980 37256 35032 37262
rect 34980 37198 35032 37204
rect 34796 37188 34848 37194
rect 34796 37130 34848 37136
rect 34520 36916 34572 36922
rect 34348 36876 34520 36904
rect 34520 36858 34572 36864
rect 34244 36168 34296 36174
rect 34244 36110 34296 36116
rect 34060 35624 34112 35630
rect 34060 35566 34112 35572
rect 34072 35086 34100 35566
rect 34060 35080 34112 35086
rect 34060 35022 34112 35028
rect 34256 33862 34284 36110
rect 34808 35894 34836 37130
rect 34992 36582 35020 37198
rect 35084 36854 35112 37334
rect 35360 37126 35388 39222
rect 35438 39200 35494 40000
rect 35990 39200 36046 40000
rect 36542 39200 36598 40000
rect 37094 39200 37150 40000
rect 37646 39200 37702 40000
rect 38198 39200 38254 40000
rect 35348 37120 35400 37126
rect 35348 37062 35400 37068
rect 35072 36848 35124 36854
rect 35072 36790 35124 36796
rect 35452 36650 35480 39200
rect 35624 37188 35676 37194
rect 35624 37130 35676 37136
rect 35440 36644 35492 36650
rect 35440 36586 35492 36592
rect 34980 36576 35032 36582
rect 34980 36518 35032 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35440 36100 35492 36106
rect 35440 36042 35492 36048
rect 34716 35866 34836 35894
rect 34610 35728 34666 35737
rect 34610 35663 34666 35672
rect 34518 35048 34574 35057
rect 34518 34983 34520 34992
rect 34572 34983 34574 34992
rect 34520 34954 34572 34960
rect 34624 34950 34652 35663
rect 34716 35494 34744 35866
rect 35348 35624 35400 35630
rect 35348 35566 35400 35572
rect 34704 35488 34756 35494
rect 34704 35430 34756 35436
rect 34612 34944 34664 34950
rect 34610 34912 34612 34921
rect 34664 34912 34666 34921
rect 34610 34847 34666 34856
rect 34518 33960 34574 33969
rect 34518 33895 34520 33904
rect 34572 33895 34574 33904
rect 34520 33866 34572 33872
rect 34244 33856 34296 33862
rect 34244 33798 34296 33804
rect 34716 31958 34744 35430
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34796 34604 34848 34610
rect 34796 34546 34848 34552
rect 34808 32026 34836 34546
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34796 32020 34848 32026
rect 34796 31962 34848 31968
rect 34704 31952 34756 31958
rect 34704 31894 34756 31900
rect 34612 31272 34664 31278
rect 34612 31214 34664 31220
rect 34520 28144 34572 28150
rect 34520 28086 34572 28092
rect 34060 26988 34112 26994
rect 34060 26930 34112 26936
rect 34072 25498 34100 26930
rect 34060 25492 34112 25498
rect 34060 25434 34112 25440
rect 34532 24750 34560 28086
rect 34624 27985 34652 31214
rect 34610 27976 34666 27985
rect 34610 27911 34666 27920
rect 34612 25696 34664 25702
rect 34612 25638 34664 25644
rect 34520 24744 34572 24750
rect 34520 24686 34572 24692
rect 34336 24608 34388 24614
rect 34336 24550 34388 24556
rect 34152 24268 34204 24274
rect 34152 24210 34204 24216
rect 34164 24070 34192 24210
rect 34348 24206 34376 24550
rect 34336 24200 34388 24206
rect 34336 24142 34388 24148
rect 34520 24200 34572 24206
rect 34520 24142 34572 24148
rect 34152 24064 34204 24070
rect 34152 24006 34204 24012
rect 34164 23662 34192 24006
rect 34532 23730 34560 24142
rect 34624 24138 34652 25638
rect 34716 25378 34744 31894
rect 34808 31414 34836 31962
rect 35256 31680 35308 31686
rect 35256 31622 35308 31628
rect 34888 31476 34940 31482
rect 34888 31418 34940 31424
rect 34796 31408 34848 31414
rect 34796 31350 34848 31356
rect 34900 31124 34928 31418
rect 35268 31346 35296 31622
rect 35256 31340 35308 31346
rect 35256 31282 35308 31288
rect 34808 31096 34928 31124
rect 34808 25702 34836 31096
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35360 27130 35388 35566
rect 35452 31090 35480 36042
rect 35636 31482 35664 37130
rect 35900 36780 35952 36786
rect 35900 36722 35952 36728
rect 35912 36650 35940 36722
rect 35900 36644 35952 36650
rect 35900 36586 35952 36592
rect 36004 35834 36032 39200
rect 36084 37256 36136 37262
rect 36084 37198 36136 37204
rect 36096 36650 36124 37198
rect 36452 36780 36504 36786
rect 36452 36722 36504 36728
rect 36084 36644 36136 36650
rect 36084 36586 36136 36592
rect 36096 36106 36124 36586
rect 36084 36100 36136 36106
rect 36084 36042 36136 36048
rect 35992 35828 36044 35834
rect 35992 35770 36044 35776
rect 35900 35488 35952 35494
rect 35900 35430 35952 35436
rect 35912 34082 35940 35430
rect 36096 35086 36124 36042
rect 36176 35692 36228 35698
rect 36176 35634 36228 35640
rect 36084 35080 36136 35086
rect 36084 35022 36136 35028
rect 35992 34536 36044 34542
rect 35992 34478 36044 34484
rect 36004 34202 36032 34478
rect 35992 34196 36044 34202
rect 35992 34138 36044 34144
rect 35912 34054 36032 34082
rect 35900 33992 35952 33998
rect 35900 33934 35952 33940
rect 35912 33454 35940 33934
rect 35900 33448 35952 33454
rect 35900 33390 35952 33396
rect 35912 32230 35940 33390
rect 35900 32224 35952 32230
rect 35900 32166 35952 32172
rect 35912 31890 35940 32166
rect 35900 31884 35952 31890
rect 35900 31826 35952 31832
rect 35624 31476 35676 31482
rect 35624 31418 35676 31424
rect 35452 31062 35848 31090
rect 35716 30660 35768 30666
rect 35716 30602 35768 30608
rect 35440 29572 35492 29578
rect 35440 29514 35492 29520
rect 35348 27124 35400 27130
rect 35348 27066 35400 27072
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35348 26376 35400 26382
rect 35348 26318 35400 26324
rect 34796 25696 34848 25702
rect 34796 25638 34848 25644
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35360 25498 35388 26318
rect 35348 25492 35400 25498
rect 35348 25434 35400 25440
rect 34716 25350 34836 25378
rect 34704 25288 34756 25294
rect 34704 25230 34756 25236
rect 34612 24132 34664 24138
rect 34612 24074 34664 24080
rect 34520 23724 34572 23730
rect 34520 23666 34572 23672
rect 34152 23656 34204 23662
rect 34152 23598 34204 23604
rect 34164 23186 34192 23598
rect 34532 23186 34560 23666
rect 34716 23322 34744 25230
rect 34808 24290 34836 25350
rect 35348 24812 35400 24818
rect 35348 24754 35400 24760
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34808 24262 34928 24290
rect 34796 24200 34848 24206
rect 34796 24142 34848 24148
rect 34808 23866 34836 24142
rect 34796 23860 34848 23866
rect 34796 23802 34848 23808
rect 34900 23610 34928 24262
rect 34808 23582 34928 23610
rect 34704 23316 34756 23322
rect 34704 23258 34756 23264
rect 34152 23180 34204 23186
rect 34152 23122 34204 23128
rect 34520 23180 34572 23186
rect 34520 23122 34572 23128
rect 34704 22636 34756 22642
rect 34704 22578 34756 22584
rect 34612 22432 34664 22438
rect 34612 22374 34664 22380
rect 34624 22030 34652 22374
rect 34716 22234 34744 22578
rect 34704 22228 34756 22234
rect 34704 22170 34756 22176
rect 34612 22024 34664 22030
rect 34612 21966 34664 21972
rect 34808 21690 34836 23582
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35360 23254 35388 24754
rect 35452 24410 35480 29514
rect 35624 27124 35676 27130
rect 35624 27066 35676 27072
rect 35532 26240 35584 26246
rect 35532 26182 35584 26188
rect 35544 26042 35572 26182
rect 35532 26036 35584 26042
rect 35532 25978 35584 25984
rect 35532 25288 35584 25294
rect 35532 25230 35584 25236
rect 35440 24404 35492 24410
rect 35440 24346 35492 24352
rect 35348 23248 35400 23254
rect 35348 23190 35400 23196
rect 34888 23112 34940 23118
rect 34888 23054 34940 23060
rect 34900 22778 34928 23054
rect 34888 22772 34940 22778
rect 34888 22714 34940 22720
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35440 21888 35492 21894
rect 35440 21830 35492 21836
rect 34796 21684 34848 21690
rect 34796 21626 34848 21632
rect 35452 21350 35480 21830
rect 35440 21344 35492 21350
rect 35440 21286 35492 21292
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34612 18216 34664 18222
rect 34612 18158 34664 18164
rect 34624 17882 34652 18158
rect 34796 18080 34848 18086
rect 34796 18022 34848 18028
rect 34612 17876 34664 17882
rect 34612 17818 34664 17824
rect 34624 17542 34652 17818
rect 34612 17536 34664 17542
rect 34612 17478 34664 17484
rect 33968 17332 34020 17338
rect 33968 17274 34020 17280
rect 34612 14272 34664 14278
rect 34612 14214 34664 14220
rect 33784 12980 33836 12986
rect 33784 12922 33836 12928
rect 33692 11008 33744 11014
rect 33692 10950 33744 10956
rect 34244 11008 34296 11014
rect 34244 10950 34296 10956
rect 33784 10668 33836 10674
rect 33784 10610 33836 10616
rect 33796 10062 33824 10610
rect 33784 10056 33836 10062
rect 33784 9998 33836 10004
rect 33600 9104 33652 9110
rect 33600 9046 33652 9052
rect 33692 6248 33744 6254
rect 33692 6190 33744 6196
rect 33600 5296 33652 5302
rect 33600 5238 33652 5244
rect 33612 3738 33640 5238
rect 33704 4826 33732 6190
rect 33796 5302 33824 9998
rect 34152 8900 34204 8906
rect 34152 8842 34204 8848
rect 34060 8832 34112 8838
rect 34060 8774 34112 8780
rect 33968 8084 34020 8090
rect 33968 8026 34020 8032
rect 33980 7410 34008 8026
rect 34072 7426 34100 8774
rect 34164 8634 34192 8842
rect 34152 8628 34204 8634
rect 34152 8570 34204 8576
rect 33968 7404 34020 7410
rect 34072 7398 34192 7426
rect 33968 7346 34020 7352
rect 34060 7268 34112 7274
rect 34060 7210 34112 7216
rect 33968 6792 34020 6798
rect 33968 6734 34020 6740
rect 33980 6458 34008 6734
rect 33968 6452 34020 6458
rect 33968 6394 34020 6400
rect 33968 6316 34020 6322
rect 33968 6258 34020 6264
rect 33784 5296 33836 5302
rect 33784 5238 33836 5244
rect 33692 4820 33744 4826
rect 33692 4762 33744 4768
rect 33600 3732 33652 3738
rect 33600 3674 33652 3680
rect 33796 3534 33824 5238
rect 33876 4616 33928 4622
rect 33876 4558 33928 4564
rect 33784 3528 33836 3534
rect 33784 3470 33836 3476
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 33784 3392 33836 3398
rect 33784 3334 33836 3340
rect 33506 3088 33562 3097
rect 33506 3023 33562 3032
rect 33520 2854 33548 3023
rect 33508 2848 33560 2854
rect 33508 2790 33560 2796
rect 33612 2650 33640 3334
rect 33796 3194 33824 3334
rect 33784 3188 33836 3194
rect 33784 3130 33836 3136
rect 33888 2774 33916 4558
rect 33980 3194 34008 6258
rect 34072 4622 34100 7210
rect 34060 4616 34112 4622
rect 34060 4558 34112 4564
rect 33968 3188 34020 3194
rect 33968 3130 34020 3136
rect 34164 3058 34192 7398
rect 34152 3052 34204 3058
rect 34152 2994 34204 3000
rect 33796 2746 33916 2774
rect 33600 2644 33652 2650
rect 33600 2586 33652 2592
rect 33796 800 33824 2746
rect 34256 2446 34284 10950
rect 34336 9104 34388 9110
rect 34336 9046 34388 9052
rect 34348 6866 34376 9046
rect 34624 8566 34652 14214
rect 34808 12850 34836 18022
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34796 12844 34848 12850
rect 34796 12786 34848 12792
rect 35348 12844 35400 12850
rect 35348 12786 35400 12792
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35360 12238 35388 12786
rect 35348 12232 35400 12238
rect 35348 12174 35400 12180
rect 35360 11762 35388 12174
rect 35348 11756 35400 11762
rect 35348 11698 35400 11704
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34796 9512 34848 9518
rect 34796 9454 34848 9460
rect 34808 9178 34836 9454
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34796 9172 34848 9178
rect 34796 9114 34848 9120
rect 34704 8968 34756 8974
rect 34704 8910 34756 8916
rect 34612 8560 34664 8566
rect 34612 8502 34664 8508
rect 34428 8492 34480 8498
rect 34428 8434 34480 8440
rect 34336 6860 34388 6866
rect 34336 6802 34388 6808
rect 34348 6458 34376 6802
rect 34440 6662 34468 8434
rect 34716 8090 34744 8910
rect 35452 8634 35480 21286
rect 35544 21146 35572 25230
rect 35636 22030 35664 27066
rect 35728 25430 35756 30602
rect 35716 25424 35768 25430
rect 35716 25366 35768 25372
rect 35716 25288 35768 25294
rect 35716 25230 35768 25236
rect 35728 24342 35756 25230
rect 35716 24336 35768 24342
rect 35716 24278 35768 24284
rect 35716 24200 35768 24206
rect 35716 24142 35768 24148
rect 35728 23322 35756 24142
rect 35820 23338 35848 31062
rect 35912 30734 35940 31826
rect 35900 30728 35952 30734
rect 35900 30670 35952 30676
rect 35900 30184 35952 30190
rect 35900 30126 35952 30132
rect 35912 29646 35940 30126
rect 35900 29640 35952 29646
rect 35900 29582 35952 29588
rect 35912 28014 35940 29582
rect 35900 28008 35952 28014
rect 35900 27950 35952 27956
rect 36004 25378 36032 34054
rect 36096 33998 36124 35022
rect 36084 33992 36136 33998
rect 36084 33934 36136 33940
rect 36084 31136 36136 31142
rect 36084 31078 36136 31084
rect 36096 25809 36124 31078
rect 36188 29850 36216 35634
rect 36266 34504 36322 34513
rect 36266 34439 36268 34448
rect 36320 34439 36322 34448
rect 36268 34410 36320 34416
rect 36280 32570 36308 34410
rect 36360 34400 36412 34406
rect 36360 34342 36412 34348
rect 36372 33522 36400 34342
rect 36360 33516 36412 33522
rect 36360 33458 36412 33464
rect 36268 32564 36320 32570
rect 36268 32506 36320 32512
rect 36464 30938 36492 36722
rect 36556 36378 36584 39200
rect 36728 37120 36780 37126
rect 36728 37062 36780 37068
rect 36544 36372 36596 36378
rect 36544 36314 36596 36320
rect 36544 36032 36596 36038
rect 36542 36000 36544 36009
rect 36596 36000 36598 36009
rect 36542 35935 36598 35944
rect 36740 35698 36768 37062
rect 37108 36310 37136 39200
rect 37096 36304 37148 36310
rect 37096 36246 37148 36252
rect 37660 35834 37688 39200
rect 38108 36780 38160 36786
rect 38108 36722 38160 36728
rect 37924 36576 37976 36582
rect 37924 36518 37976 36524
rect 37740 36168 37792 36174
rect 37740 36110 37792 36116
rect 37648 35828 37700 35834
rect 37648 35770 37700 35776
rect 36728 35692 36780 35698
rect 36728 35634 36780 35640
rect 37648 35692 37700 35698
rect 37648 35634 37700 35640
rect 37660 34950 37688 35634
rect 36728 34944 36780 34950
rect 36728 34886 36780 34892
rect 37648 34944 37700 34950
rect 37648 34886 37700 34892
rect 36452 30932 36504 30938
rect 36452 30874 36504 30880
rect 36176 29844 36228 29850
rect 36176 29786 36228 29792
rect 36188 29730 36216 29786
rect 36188 29702 36308 29730
rect 36176 28484 36228 28490
rect 36176 28426 36228 28432
rect 36082 25800 36138 25809
rect 36082 25735 36138 25744
rect 36004 25350 36124 25378
rect 35992 25220 36044 25226
rect 35992 25162 36044 25168
rect 36004 24682 36032 25162
rect 35992 24676 36044 24682
rect 35992 24618 36044 24624
rect 35820 23322 35940 23338
rect 35716 23316 35768 23322
rect 35820 23316 35952 23322
rect 35820 23310 35900 23316
rect 35716 23258 35768 23264
rect 35900 23258 35952 23264
rect 35900 22976 35952 22982
rect 35900 22918 35952 22924
rect 35716 22704 35768 22710
rect 35716 22646 35768 22652
rect 35624 22024 35676 22030
rect 35624 21966 35676 21972
rect 35532 21140 35584 21146
rect 35532 21082 35584 21088
rect 35728 16574 35756 22646
rect 35808 22568 35860 22574
rect 35808 22510 35860 22516
rect 35820 22098 35848 22510
rect 35912 22234 35940 22918
rect 35900 22228 35952 22234
rect 35900 22170 35952 22176
rect 35808 22092 35860 22098
rect 35808 22034 35860 22040
rect 35820 21010 35848 22034
rect 35900 21072 35952 21078
rect 35900 21014 35952 21020
rect 35808 21004 35860 21010
rect 35808 20946 35860 20952
rect 35808 20868 35860 20874
rect 35808 20810 35860 20816
rect 35636 16546 35756 16574
rect 35532 11144 35584 11150
rect 35532 11086 35584 11092
rect 35544 10742 35572 11086
rect 35532 10736 35584 10742
rect 35532 10678 35584 10684
rect 35544 9654 35572 10678
rect 35532 9648 35584 9654
rect 35532 9590 35584 9596
rect 35544 8974 35572 9590
rect 35636 9382 35664 16546
rect 35624 9376 35676 9382
rect 35624 9318 35676 9324
rect 35532 8968 35584 8974
rect 35532 8910 35584 8916
rect 35440 8628 35492 8634
rect 35440 8570 35492 8576
rect 35348 8288 35400 8294
rect 35348 8230 35400 8236
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34704 8084 34756 8090
rect 34704 8026 34756 8032
rect 35360 7954 35388 8230
rect 35348 7948 35400 7954
rect 35348 7890 35400 7896
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 34808 7546 34836 7822
rect 34796 7540 34848 7546
rect 34796 7482 34848 7488
rect 35360 7206 35388 7890
rect 35348 7200 35400 7206
rect 35348 7142 35400 7148
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35360 6866 35388 7142
rect 35348 6860 35400 6866
rect 35348 6802 35400 6808
rect 34428 6656 34480 6662
rect 34428 6598 34480 6604
rect 34336 6452 34388 6458
rect 34336 6394 34388 6400
rect 34704 6316 34756 6322
rect 34704 6258 34756 6264
rect 34716 5914 34744 6258
rect 35360 6118 35388 6802
rect 34796 6112 34848 6118
rect 34796 6054 34848 6060
rect 35348 6112 35400 6118
rect 35348 6054 35400 6060
rect 34704 5908 34756 5914
rect 34704 5850 34756 5856
rect 34808 5642 34836 6054
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35360 5778 35388 6054
rect 35348 5772 35400 5778
rect 35348 5714 35400 5720
rect 34796 5636 34848 5642
rect 34796 5578 34848 5584
rect 34520 5568 34572 5574
rect 34520 5510 34572 5516
rect 34532 4826 34560 5510
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34520 4820 34572 4826
rect 34520 4762 34572 4768
rect 35360 4758 35388 5714
rect 35348 4752 35400 4758
rect 35348 4694 35400 4700
rect 35452 4690 35480 8570
rect 35636 8022 35664 9318
rect 35820 8566 35848 20810
rect 35912 19922 35940 21014
rect 35900 19916 35952 19922
rect 35900 19858 35952 19864
rect 35912 19378 35940 19858
rect 36096 19514 36124 25350
rect 36188 24682 36216 28426
rect 36176 24676 36228 24682
rect 36176 24618 36228 24624
rect 36280 22030 36308 29702
rect 36360 25696 36412 25702
rect 36360 25638 36412 25644
rect 36372 25362 36400 25638
rect 36360 25356 36412 25362
rect 36360 25298 36412 25304
rect 36464 24290 36492 30874
rect 36544 29572 36596 29578
rect 36544 29514 36596 29520
rect 36556 24410 36584 29514
rect 36636 26580 36688 26586
rect 36636 26522 36688 26528
rect 36648 25702 36676 26522
rect 36740 26042 36768 34886
rect 37096 33924 37148 33930
rect 37096 33866 37148 33872
rect 36820 28552 36872 28558
rect 36872 28500 37044 28506
rect 36820 28494 37044 28500
rect 36832 28478 37044 28494
rect 37016 28014 37044 28478
rect 37004 28008 37056 28014
rect 37004 27950 37056 27956
rect 37016 27470 37044 27950
rect 37004 27464 37056 27470
rect 37004 27406 37056 27412
rect 37016 26586 37044 27406
rect 37004 26580 37056 26586
rect 37004 26522 37056 26528
rect 37108 26234 37136 33866
rect 36924 26206 37136 26234
rect 36728 26036 36780 26042
rect 36728 25978 36780 25984
rect 36636 25696 36688 25702
rect 36636 25638 36688 25644
rect 36544 24404 36596 24410
rect 36544 24346 36596 24352
rect 36372 24262 36492 24290
rect 36372 22778 36400 24262
rect 36452 24200 36504 24206
rect 36452 24142 36504 24148
rect 36360 22772 36412 22778
rect 36360 22714 36412 22720
rect 36268 22024 36320 22030
rect 36268 21966 36320 21972
rect 36268 21548 36320 21554
rect 36268 21490 36320 21496
rect 36280 20058 36308 21490
rect 36464 21486 36492 24142
rect 36452 21480 36504 21486
rect 36452 21422 36504 21428
rect 36740 21146 36768 25978
rect 36820 24744 36872 24750
rect 36820 24686 36872 24692
rect 36832 24614 36860 24686
rect 36820 24608 36872 24614
rect 36820 24550 36872 24556
rect 36728 21140 36780 21146
rect 36728 21082 36780 21088
rect 36740 20942 36768 21082
rect 36832 21078 36860 24550
rect 36924 22817 36952 26206
rect 37660 24954 37688 34886
rect 37752 33658 37780 36110
rect 37936 35894 37964 36518
rect 37936 35866 38056 35894
rect 37832 35012 37884 35018
rect 37832 34954 37884 34960
rect 37740 33652 37792 33658
rect 37740 33594 37792 33600
rect 37844 26042 37872 34954
rect 37924 29844 37976 29850
rect 37924 29786 37976 29792
rect 37832 26036 37884 26042
rect 37832 25978 37884 25984
rect 37936 25242 37964 29786
rect 38028 28762 38056 35866
rect 38120 29850 38148 36722
rect 38212 34610 38240 39200
rect 38292 37120 38344 37126
rect 38292 37062 38344 37068
rect 38200 34604 38252 34610
rect 38200 34546 38252 34552
rect 38108 29844 38160 29850
rect 38108 29786 38160 29792
rect 38016 28756 38068 28762
rect 38016 28698 38068 28704
rect 38028 26234 38056 28698
rect 38304 26234 38332 37062
rect 38028 26206 38148 26234
rect 38016 25900 38068 25906
rect 38016 25842 38068 25848
rect 37752 25214 37964 25242
rect 37648 24948 37700 24954
rect 37648 24890 37700 24896
rect 37752 23798 37780 25214
rect 37832 25152 37884 25158
rect 37832 25094 37884 25100
rect 37844 24682 37872 25094
rect 37832 24676 37884 24682
rect 37832 24618 37884 24624
rect 37924 24608 37976 24614
rect 37924 24550 37976 24556
rect 37936 24206 37964 24550
rect 38028 24410 38056 25842
rect 38016 24404 38068 24410
rect 38016 24346 38068 24352
rect 37924 24200 37976 24206
rect 37924 24142 37976 24148
rect 37740 23792 37792 23798
rect 37740 23734 37792 23740
rect 37096 23520 37148 23526
rect 37096 23462 37148 23468
rect 37004 23112 37056 23118
rect 37004 23054 37056 23060
rect 36910 22808 36966 22817
rect 36910 22743 36966 22752
rect 37016 21690 37044 23054
rect 37004 21684 37056 21690
rect 37004 21626 37056 21632
rect 36820 21072 36872 21078
rect 36820 21014 36872 21020
rect 36728 20936 36780 20942
rect 36728 20878 36780 20884
rect 36268 20052 36320 20058
rect 36268 19994 36320 20000
rect 36450 19952 36506 19961
rect 36450 19887 36506 19896
rect 36464 19854 36492 19887
rect 36452 19848 36504 19854
rect 36452 19790 36504 19796
rect 36084 19508 36136 19514
rect 36084 19450 36136 19456
rect 35900 19372 35952 19378
rect 35900 19314 35952 19320
rect 36096 18970 36124 19450
rect 36544 19304 36596 19310
rect 36544 19246 36596 19252
rect 36084 18964 36136 18970
rect 36084 18906 36136 18912
rect 36268 15564 36320 15570
rect 36268 15506 36320 15512
rect 36280 14482 36308 15506
rect 36452 15360 36504 15366
rect 36452 15302 36504 15308
rect 36268 14476 36320 14482
rect 36268 14418 36320 14424
rect 36464 13938 36492 15302
rect 36556 14482 36584 19246
rect 36912 15360 36964 15366
rect 36912 15302 36964 15308
rect 36544 14476 36596 14482
rect 36596 14436 36676 14464
rect 36544 14418 36596 14424
rect 36544 14272 36596 14278
rect 36544 14214 36596 14220
rect 36452 13932 36504 13938
rect 36452 13874 36504 13880
rect 36268 13728 36320 13734
rect 36268 13670 36320 13676
rect 36280 12434 36308 13670
rect 36280 12406 36400 12434
rect 36372 12170 36400 12406
rect 36360 12164 36412 12170
rect 36360 12106 36412 12112
rect 35808 8560 35860 8566
rect 35808 8502 35860 8508
rect 35624 8016 35676 8022
rect 35624 7958 35676 7964
rect 35820 7834 35848 8502
rect 35728 7806 35848 7834
rect 36176 7880 36228 7886
rect 36176 7822 36228 7828
rect 35440 4684 35492 4690
rect 35440 4626 35492 4632
rect 35072 4480 35124 4486
rect 35072 4422 35124 4428
rect 35084 4282 35112 4422
rect 35452 4282 35480 4626
rect 35072 4276 35124 4282
rect 35072 4218 35124 4224
rect 35440 4276 35492 4282
rect 35440 4218 35492 4224
rect 35728 4078 35756 7806
rect 35808 7744 35860 7750
rect 35808 7686 35860 7692
rect 35716 4072 35768 4078
rect 35716 4014 35768 4020
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35348 3528 35400 3534
rect 35348 3470 35400 3476
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 34336 2848 34388 2854
rect 34336 2790 34388 2796
rect 34244 2440 34296 2446
rect 34244 2382 34296 2388
rect 34348 800 34376 2790
rect 34808 2446 34836 3334
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 34900 870 35020 898
rect 34900 800 34928 870
rect 27816 734 28120 762
rect 28262 0 28318 800
rect 28814 0 28870 800
rect 29366 0 29422 800
rect 29918 0 29974 800
rect 30470 0 30526 800
rect 31022 0 31078 800
rect 31574 0 31630 800
rect 32126 0 32182 800
rect 32678 0 32734 800
rect 33230 0 33286 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34886 0 34942 800
rect 34992 762 35020 870
rect 35360 762 35388 3470
rect 35728 3194 35756 4014
rect 35820 3398 35848 7686
rect 35992 7404 36044 7410
rect 35992 7346 36044 7352
rect 35900 7268 35952 7274
rect 35900 7210 35952 7216
rect 35912 5710 35940 7210
rect 36004 5914 36032 7346
rect 36188 6866 36216 7822
rect 36176 6860 36228 6866
rect 36176 6802 36228 6808
rect 36084 6656 36136 6662
rect 36084 6598 36136 6604
rect 35992 5908 36044 5914
rect 35992 5850 36044 5856
rect 35900 5704 35952 5710
rect 35900 5646 35952 5652
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 35716 3188 35768 3194
rect 35716 3130 35768 3136
rect 35912 2774 35940 5646
rect 36096 4842 36124 6598
rect 36188 5846 36216 6802
rect 36176 5840 36228 5846
rect 36176 5782 36228 5788
rect 36188 5302 36216 5782
rect 36176 5296 36228 5302
rect 36176 5238 36228 5244
rect 36004 4814 36124 4842
rect 36004 4146 36032 4814
rect 36188 4706 36216 5238
rect 36452 5092 36504 5098
rect 36452 5034 36504 5040
rect 36268 5024 36320 5030
rect 36268 4966 36320 4972
rect 36096 4678 36216 4706
rect 36096 4622 36124 4678
rect 36280 4622 36308 4966
rect 36084 4616 36136 4622
rect 36084 4558 36136 4564
rect 36268 4616 36320 4622
rect 36268 4558 36320 4564
rect 36096 4214 36124 4558
rect 36084 4208 36136 4214
rect 36084 4150 36136 4156
rect 36360 4208 36412 4214
rect 36360 4150 36412 4156
rect 35992 4140 36044 4146
rect 35992 4082 36044 4088
rect 36372 3602 36400 4150
rect 36464 4146 36492 5034
rect 36556 4554 36584 14214
rect 36648 13530 36676 14436
rect 36636 13524 36688 13530
rect 36636 13466 36688 13472
rect 36636 6112 36688 6118
rect 36636 6054 36688 6060
rect 36544 4548 36596 4554
rect 36544 4490 36596 4496
rect 36452 4140 36504 4146
rect 36452 4082 36504 4088
rect 36544 3664 36596 3670
rect 36544 3606 36596 3612
rect 36360 3596 36412 3602
rect 36360 3538 36412 3544
rect 35990 3496 36046 3505
rect 35990 3431 35992 3440
rect 36044 3431 36046 3440
rect 35992 3402 36044 3408
rect 35992 3188 36044 3194
rect 35992 3130 36044 3136
rect 35820 2746 35940 2774
rect 35452 870 35572 898
rect 35452 800 35480 870
rect 34992 734 35388 762
rect 35438 0 35494 800
rect 35544 762 35572 870
rect 35820 762 35848 2746
rect 36004 800 36032 3130
rect 36372 3058 36400 3538
rect 36360 3052 36412 3058
rect 36360 2994 36412 3000
rect 36372 2774 36400 2994
rect 36372 2746 36492 2774
rect 36464 2650 36492 2746
rect 36452 2644 36504 2650
rect 36452 2586 36504 2592
rect 36556 800 36584 3606
rect 36648 2446 36676 6054
rect 36924 5370 36952 15302
rect 37004 8832 37056 8838
rect 37004 8774 37056 8780
rect 36912 5364 36964 5370
rect 36912 5306 36964 5312
rect 37016 3534 37044 8774
rect 37108 8090 37136 23462
rect 38120 22438 38148 26206
rect 38212 26206 38332 26234
rect 38212 25158 38240 26206
rect 38200 25152 38252 25158
rect 38200 25094 38252 25100
rect 38108 22432 38160 22438
rect 38108 22374 38160 22380
rect 37372 21888 37424 21894
rect 37372 21830 37424 21836
rect 37384 16574 37412 21830
rect 37464 19712 37516 19718
rect 37464 19654 37516 19660
rect 37292 16546 37412 16574
rect 37292 14362 37320 16546
rect 37476 15450 37504 19654
rect 37740 17536 37792 17542
rect 37740 17478 37792 17484
rect 37752 16574 37780 17478
rect 37384 15422 37504 15450
rect 37568 16546 37780 16574
rect 37384 15366 37412 15422
rect 37372 15360 37424 15366
rect 37372 15302 37424 15308
rect 37200 14334 37320 14362
rect 37200 12730 37228 14334
rect 37280 14272 37332 14278
rect 37280 14214 37332 14220
rect 37292 12850 37320 14214
rect 37280 12844 37332 12850
rect 37280 12786 37332 12792
rect 37200 12702 37320 12730
rect 37096 8084 37148 8090
rect 37096 8026 37148 8032
rect 37108 7546 37136 8026
rect 37096 7540 37148 7546
rect 37096 7482 37148 7488
rect 37292 7478 37320 12702
rect 37384 12442 37412 15302
rect 37464 13252 37516 13258
rect 37464 13194 37516 13200
rect 37476 12986 37504 13194
rect 37464 12980 37516 12986
rect 37464 12922 37516 12928
rect 37372 12436 37424 12442
rect 37372 12378 37424 12384
rect 37370 8392 37426 8401
rect 37370 8327 37372 8336
rect 37424 8327 37426 8336
rect 37372 8298 37424 8304
rect 37280 7472 37332 7478
rect 37280 7414 37332 7420
rect 37188 6792 37240 6798
rect 37188 6734 37240 6740
rect 37200 4010 37228 6734
rect 37292 5896 37320 7414
rect 37384 6066 37412 8298
rect 37568 6769 37596 16546
rect 37924 15360 37976 15366
rect 37924 15302 37976 15308
rect 37936 12434 37964 15302
rect 38108 13320 38160 13326
rect 38108 13262 38160 13268
rect 37844 12406 37964 12434
rect 37844 11082 37872 12406
rect 38120 12238 38148 13262
rect 38108 12232 38160 12238
rect 38108 12174 38160 12180
rect 38120 11218 38148 12174
rect 38108 11212 38160 11218
rect 38108 11154 38160 11160
rect 37832 11076 37884 11082
rect 37832 11018 37884 11024
rect 38016 10464 38068 10470
rect 38016 10406 38068 10412
rect 37648 9920 37700 9926
rect 37648 9862 37700 9868
rect 37832 9920 37884 9926
rect 37832 9862 37884 9868
rect 37554 6760 37610 6769
rect 37476 6718 37554 6746
rect 37476 6225 37504 6718
rect 37554 6695 37610 6704
rect 37556 6656 37608 6662
rect 37556 6598 37608 6604
rect 37462 6216 37518 6225
rect 37568 6186 37596 6598
rect 37462 6151 37518 6160
rect 37556 6180 37608 6186
rect 37556 6122 37608 6128
rect 37384 6038 37596 6066
rect 37372 5908 37424 5914
rect 37292 5868 37372 5896
rect 37372 5850 37424 5856
rect 37372 5296 37424 5302
rect 37372 5238 37424 5244
rect 37384 4758 37412 5238
rect 37464 5228 37516 5234
rect 37464 5170 37516 5176
rect 37476 4826 37504 5170
rect 37464 4820 37516 4826
rect 37464 4762 37516 4768
rect 37372 4752 37424 4758
rect 37372 4694 37424 4700
rect 37188 4004 37240 4010
rect 37188 3946 37240 3952
rect 37280 3936 37332 3942
rect 37280 3878 37332 3884
rect 37004 3528 37056 3534
rect 37002 3496 37004 3505
rect 37056 3496 37058 3505
rect 37002 3431 37058 3440
rect 37292 3126 37320 3878
rect 37568 3466 37596 6038
rect 37660 3534 37688 9862
rect 37740 9376 37792 9382
rect 37740 9318 37792 9324
rect 37752 4146 37780 9318
rect 37740 4140 37792 4146
rect 37740 4082 37792 4088
rect 37752 3602 37780 4082
rect 37740 3596 37792 3602
rect 37740 3538 37792 3544
rect 37648 3528 37700 3534
rect 37648 3470 37700 3476
rect 37556 3460 37608 3466
rect 37556 3402 37608 3408
rect 37660 3210 37688 3470
rect 37568 3182 37688 3210
rect 37280 3120 37332 3126
rect 37280 3062 37332 3068
rect 37568 2854 37596 3182
rect 37648 3120 37700 3126
rect 37648 3062 37700 3068
rect 37556 2848 37608 2854
rect 37556 2790 37608 2796
rect 37554 2544 37610 2553
rect 37554 2479 37556 2488
rect 37608 2479 37610 2488
rect 37556 2450 37608 2456
rect 36636 2440 36688 2446
rect 36636 2382 36688 2388
rect 37096 2440 37148 2446
rect 37096 2382 37148 2388
rect 37108 800 37136 2382
rect 37660 800 37688 3062
rect 37844 2446 37872 9862
rect 37924 8832 37976 8838
rect 37924 8774 37976 8780
rect 37936 4622 37964 8774
rect 37924 4616 37976 4622
rect 37924 4558 37976 4564
rect 37936 3194 37964 4558
rect 37924 3188 37976 3194
rect 37924 3130 37976 3136
rect 38028 3126 38056 10406
rect 38108 8356 38160 8362
rect 38108 8298 38160 8304
rect 38120 5234 38148 8298
rect 38200 7880 38252 7886
rect 38200 7822 38252 7828
rect 38108 5228 38160 5234
rect 38108 5170 38160 5176
rect 38120 3670 38148 5170
rect 38108 3664 38160 3670
rect 38108 3606 38160 3612
rect 38016 3120 38068 3126
rect 38016 3062 38068 3068
rect 37832 2440 37884 2446
rect 37832 2382 37884 2388
rect 38212 800 38240 7822
rect 38290 6760 38346 6769
rect 38290 6695 38346 6704
rect 38304 2854 38332 6695
rect 38292 2848 38344 2854
rect 38292 2790 38344 2796
rect 35544 734 35848 762
rect 35990 0 36046 800
rect 36542 0 36598 800
rect 37094 0 37150 800
rect 37646 0 37702 800
rect 38198 0 38254 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 10230 36080 10286 36136
rect 8850 25200 8906 25256
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 9494 27376 9550 27432
rect 9954 28056 10010 28112
rect 10230 26852 10286 26888
rect 10230 26832 10232 26852
rect 10232 26832 10284 26852
rect 10284 26832 10286 26852
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4986 2352 5042 2408
rect 5170 2896 5226 2952
rect 6182 3612 6184 3632
rect 6184 3612 6236 3632
rect 6236 3612 6238 3632
rect 6182 3576 6238 3612
rect 7194 3712 7250 3768
rect 10230 25372 10232 25392
rect 10232 25372 10284 25392
rect 10284 25372 10286 25392
rect 10230 25336 10286 25372
rect 10230 8880 10286 8936
rect 9678 5616 9734 5672
rect 9402 3884 9404 3904
rect 9404 3884 9456 3904
rect 9456 3884 9458 3904
rect 9402 3848 9458 3884
rect 9126 3576 9182 3632
rect 12438 35264 12494 35320
rect 12070 34584 12126 34640
rect 12254 34176 12310 34232
rect 12346 29028 12402 29064
rect 12346 29008 12348 29028
rect 12348 29008 12400 29028
rect 12400 29008 12402 29028
rect 12346 28484 12402 28520
rect 12346 28464 12348 28484
rect 12348 28464 12400 28484
rect 12400 28464 12402 28484
rect 11886 26288 11942 26344
rect 10874 10104 10930 10160
rect 11702 10532 11758 10568
rect 11702 10512 11704 10532
rect 11704 10512 11756 10532
rect 11756 10512 11758 10532
rect 13266 32272 13322 32328
rect 13174 29144 13230 29200
rect 10506 5208 10562 5264
rect 11058 5752 11114 5808
rect 10414 3712 10470 3768
rect 9954 3168 10010 3224
rect 9954 2644 10010 2680
rect 9954 2624 9956 2644
rect 9956 2624 10008 2644
rect 10008 2624 10010 2644
rect 9310 1944 9366 2000
rect 10598 4004 10654 4040
rect 10598 3984 10600 4004
rect 10600 3984 10652 4004
rect 10652 3984 10654 4004
rect 11702 6976 11758 7032
rect 11978 3576 12034 3632
rect 11518 3304 11574 3360
rect 12254 4120 12310 4176
rect 12162 3304 12218 3360
rect 12806 9460 12808 9480
rect 12808 9460 12860 9480
rect 12860 9460 12862 9480
rect 12806 9424 12862 9460
rect 13634 31728 13690 31784
rect 13542 29724 13544 29744
rect 13544 29724 13596 29744
rect 13596 29724 13598 29744
rect 13542 29688 13598 29724
rect 14830 32272 14886 32328
rect 14278 29552 14334 29608
rect 12346 3712 12402 3768
rect 12898 5908 12954 5944
rect 12898 5888 12900 5908
rect 12900 5888 12952 5908
rect 12952 5888 12954 5908
rect 12714 3984 12770 4040
rect 13358 6704 13414 6760
rect 13174 3984 13230 4040
rect 13542 3984 13598 4040
rect 13542 3576 13598 3632
rect 15290 12280 15346 12336
rect 15198 11192 15254 11248
rect 14830 9968 14886 10024
rect 13726 9016 13782 9072
rect 13726 4528 13782 4584
rect 13726 3848 13782 3904
rect 13818 2624 13874 2680
rect 13082 1808 13138 1864
rect 17682 36760 17738 36816
rect 16854 31048 16910 31104
rect 16486 30232 16542 30288
rect 16854 27940 16910 27976
rect 16854 27920 16856 27940
rect 16856 27920 16908 27940
rect 16908 27920 16910 27940
rect 16394 26968 16450 27024
rect 16210 13368 16266 13424
rect 15106 7792 15162 7848
rect 17038 25916 17040 25936
rect 17040 25916 17092 25936
rect 17092 25916 17094 25936
rect 17038 25880 17094 25916
rect 16670 25608 16726 25664
rect 16302 9968 16358 10024
rect 14738 3032 14794 3088
rect 15106 2760 15162 2816
rect 15382 4120 15438 4176
rect 16486 11600 16542 11656
rect 16670 11056 16726 11112
rect 15750 6160 15806 6216
rect 15842 5072 15898 5128
rect 16302 3168 16358 3224
rect 18326 33924 18382 33960
rect 18326 33904 18328 33924
rect 18328 33904 18380 33924
rect 18380 33904 18382 33924
rect 17682 31048 17738 31104
rect 17038 11056 17094 11112
rect 16946 9152 17002 9208
rect 16946 5752 17002 5808
rect 19062 36080 19118 36136
rect 18418 25472 18474 25528
rect 18326 17176 18382 17232
rect 17406 7384 17462 7440
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19338 35692 19394 35728
rect 19338 35672 19340 35692
rect 19340 35672 19392 35692
rect 19392 35672 19394 35692
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19982 34992 20038 35048
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19062 30232 19118 30288
rect 18694 27548 18696 27568
rect 18696 27548 18748 27568
rect 18748 27548 18750 27568
rect 18694 27512 18750 27548
rect 18694 13776 18750 13832
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19522 26444 19578 26480
rect 19522 26424 19524 26444
rect 19524 26424 19576 26444
rect 19576 26424 19578 26444
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 20074 23704 20130 23760
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 17958 11192 18014 11248
rect 17958 7268 18014 7304
rect 17958 7248 17960 7268
rect 17960 7248 18012 7268
rect 18012 7248 18014 7268
rect 17590 5752 17646 5808
rect 16670 3032 16726 3088
rect 16946 3052 17002 3088
rect 16946 3032 16948 3052
rect 16948 3032 17000 3052
rect 17000 3032 17002 3052
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 21178 36488 21234 36544
rect 21086 36352 21142 36408
rect 21730 36216 21786 36272
rect 20810 33088 20866 33144
rect 22374 36488 22430 36544
rect 22742 35808 22798 35864
rect 21638 35128 21694 35184
rect 20534 29280 20590 29336
rect 20994 29416 21050 29472
rect 20626 26424 20682 26480
rect 20442 24792 20498 24848
rect 20074 13232 20130 13288
rect 18142 4256 18198 4312
rect 18234 4120 18290 4176
rect 16946 2488 17002 2544
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19062 6296 19118 6352
rect 18694 6024 18750 6080
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 18786 2488 18842 2544
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 20258 8336 20314 8392
rect 19246 3712 19302 3768
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19706 3596 19762 3632
rect 19706 3576 19708 3596
rect 19708 3576 19760 3596
rect 19760 3576 19762 3596
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20626 14612 20682 14648
rect 20626 14592 20628 14612
rect 20628 14592 20680 14612
rect 20680 14592 20682 14612
rect 20626 12144 20682 12200
rect 20442 8508 20444 8528
rect 20444 8508 20496 8528
rect 20496 8508 20498 8528
rect 20442 8472 20498 8508
rect 19614 2896 19670 2952
rect 20534 4256 20590 4312
rect 20442 3576 20498 3632
rect 19614 2372 19670 2408
rect 19614 2352 19616 2372
rect 19616 2352 19668 2372
rect 19668 2352 19670 2372
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21454 26968 21510 27024
rect 20810 5616 20866 5672
rect 20810 3984 20866 4040
rect 20810 3576 20866 3632
rect 21086 9016 21142 9072
rect 22190 34312 22246 34368
rect 21822 29280 21878 29336
rect 21638 12280 21694 12336
rect 21730 11056 21786 11112
rect 22742 33516 22798 33552
rect 22742 33496 22744 33516
rect 22744 33496 22796 33516
rect 22796 33496 22798 33516
rect 22742 32988 22744 33008
rect 22744 32988 22796 33008
rect 22796 32988 22798 33008
rect 22742 32952 22798 32988
rect 22742 32816 22798 32872
rect 22558 25880 22614 25936
rect 24122 36896 24178 36952
rect 23386 36780 23442 36816
rect 23386 36760 23388 36780
rect 23388 36760 23440 36780
rect 23440 36760 23442 36780
rect 23386 36644 23442 36680
rect 23386 36624 23388 36644
rect 23388 36624 23440 36644
rect 23440 36624 23442 36644
rect 23386 35400 23442 35456
rect 23386 34740 23442 34776
rect 23386 34720 23388 34740
rect 23388 34720 23440 34740
rect 23440 34720 23442 34740
rect 24674 36896 24730 36952
rect 24306 35944 24362 36000
rect 24582 36080 24638 36136
rect 24122 34448 24178 34504
rect 23386 32544 23442 32600
rect 23662 25200 23718 25256
rect 21822 9968 21878 10024
rect 23386 11600 23442 11656
rect 23386 10104 23442 10160
rect 24582 34060 24638 34096
rect 25410 36624 25466 36680
rect 25134 35808 25190 35864
rect 25778 36760 25834 36816
rect 25410 35400 25466 35456
rect 24582 34040 24584 34060
rect 24584 34040 24636 34060
rect 24636 34040 24638 34060
rect 24122 33224 24178 33280
rect 24398 31728 24454 31784
rect 24398 29452 24400 29472
rect 24400 29452 24452 29472
rect 24452 29452 24454 29472
rect 24398 29416 24454 29452
rect 24674 29688 24730 29744
rect 24398 25336 24454 25392
rect 25042 29144 25098 29200
rect 24858 28056 24914 28112
rect 24858 27396 24914 27432
rect 24858 27376 24860 27396
rect 24860 27376 24912 27396
rect 24912 27376 24914 27396
rect 25226 26832 25282 26888
rect 26146 36488 26202 36544
rect 26330 36760 26386 36816
rect 26238 35808 26294 35864
rect 26974 36216 27030 36272
rect 26974 34584 27030 34640
rect 28170 36916 28226 36952
rect 28170 36896 28172 36916
rect 28172 36896 28224 36916
rect 28224 36896 28226 36916
rect 28998 35264 29054 35320
rect 27802 34176 27858 34232
rect 26330 33224 26386 33280
rect 27250 32544 27306 32600
rect 27618 29008 27674 29064
rect 26974 28464 27030 28520
rect 29182 34312 29238 34368
rect 28998 33088 29054 33144
rect 28354 31084 28356 31104
rect 28356 31084 28408 31104
rect 28408 31084 28410 31104
rect 28354 31048 28410 31084
rect 27618 26288 27674 26344
rect 27986 25472 28042 25528
rect 27710 24792 27766 24848
rect 24490 13404 24492 13424
rect 24492 13404 24544 13424
rect 24544 13404 24546 13424
rect 24490 13368 24546 13404
rect 22006 7792 22062 7848
rect 21638 6704 21694 6760
rect 22282 7248 22338 7304
rect 22374 6840 22430 6896
rect 22650 5888 22706 5944
rect 21822 5208 21878 5264
rect 22374 4548 22430 4584
rect 22374 4528 22376 4548
rect 22376 4528 22428 4548
rect 22428 4528 22430 4548
rect 21638 3848 21694 3904
rect 23570 6976 23626 7032
rect 24950 15156 25006 15192
rect 24950 15136 24952 15156
rect 24952 15136 25004 15156
rect 25004 15136 25006 15156
rect 25226 9424 25282 9480
rect 24950 9288 25006 9344
rect 24030 8880 24086 8936
rect 28906 25880 28962 25936
rect 26422 14612 26478 14648
rect 26422 14592 26424 14612
rect 26424 14592 26476 14612
rect 26476 14592 26478 14612
rect 26238 10512 26294 10568
rect 26422 9172 26478 9208
rect 26422 9152 26424 9172
rect 26424 9152 26476 9172
rect 26476 9152 26478 9172
rect 26238 8492 26294 8528
rect 26238 8472 26240 8492
rect 26240 8472 26292 8492
rect 26292 8472 26294 8492
rect 26146 6024 26202 6080
rect 24582 4120 24638 4176
rect 24582 2760 24638 2816
rect 24214 1944 24270 2000
rect 25870 3576 25926 3632
rect 25502 3440 25558 3496
rect 26422 5072 26478 5128
rect 27710 12164 27766 12200
rect 27710 12144 27712 12164
rect 27712 12144 27764 12164
rect 27764 12144 27766 12164
rect 30286 36100 30342 36136
rect 30286 36080 30288 36100
rect 30288 36080 30340 36100
rect 30340 36080 30342 36100
rect 29550 29552 29606 29608
rect 31022 32292 31078 32328
rect 31022 32272 31024 32292
rect 31024 32272 31076 32292
rect 31076 32272 31078 32292
rect 29550 13232 29606 13288
rect 29366 9324 29368 9344
rect 29368 9324 29420 9344
rect 29420 9324 29422 9344
rect 27618 5752 27674 5808
rect 28998 6316 29054 6352
rect 28998 6296 29000 6316
rect 29000 6296 29052 6316
rect 29052 6296 29054 6316
rect 29366 9288 29422 9324
rect 28078 3712 28134 3768
rect 27710 1808 27766 1864
rect 28446 4276 28502 4312
rect 28446 4256 28448 4276
rect 28448 4256 28500 4276
rect 28500 4256 28502 4276
rect 28998 3732 29054 3768
rect 28998 3712 29000 3732
rect 29000 3712 29052 3732
rect 29052 3712 29054 3732
rect 31390 35164 31392 35184
rect 31392 35164 31444 35184
rect 31444 35164 31446 35184
rect 31390 35128 31446 35164
rect 31206 26016 31262 26072
rect 30930 23704 30986 23760
rect 31850 34720 31906 34776
rect 31666 34040 31722 34096
rect 31758 27512 31814 27568
rect 33966 36352 34022 36408
rect 33046 33496 33102 33552
rect 33322 32836 33378 32872
rect 33322 32816 33324 32836
rect 33324 32816 33376 32836
rect 33376 32816 33378 32836
rect 32310 22772 32366 22808
rect 32310 22752 32312 22772
rect 32312 22752 32364 22772
rect 32364 22752 32366 22772
rect 30378 7420 30380 7440
rect 30380 7420 30432 7440
rect 30432 7420 30434 7440
rect 30378 7384 30434 7420
rect 31758 3712 31814 3768
rect 31758 1672 31814 1728
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34610 35672 34666 35728
rect 34518 35012 34574 35048
rect 34518 34992 34520 35012
rect 34520 34992 34572 35012
rect 34572 34992 34574 35012
rect 34610 34892 34612 34912
rect 34612 34892 34664 34912
rect 34664 34892 34666 34912
rect 34610 34856 34666 34892
rect 34518 33924 34574 33960
rect 34518 33904 34520 33924
rect 34520 33904 34572 33924
rect 34572 33904 34574 33924
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34610 27920 34666 27976
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 33506 3032 33562 3088
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 36266 34468 36322 34504
rect 36266 34448 36268 34468
rect 36268 34448 36320 34468
rect 36320 34448 36322 34468
rect 36542 35980 36544 36000
rect 36544 35980 36596 36000
rect 36596 35980 36598 36000
rect 36542 35944 36598 35980
rect 36082 25744 36138 25800
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 36910 22752 36966 22808
rect 36450 19896 36506 19952
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35990 3460 36046 3496
rect 35990 3440 35992 3460
rect 35992 3440 36044 3460
rect 36044 3440 36046 3460
rect 37370 8356 37426 8392
rect 37370 8336 37372 8356
rect 37372 8336 37424 8356
rect 37424 8336 37426 8356
rect 37554 6704 37610 6760
rect 37462 6160 37518 6216
rect 37002 3476 37004 3496
rect 37004 3476 37056 3496
rect 37056 3476 37058 3496
rect 37002 3440 37058 3476
rect 37554 2508 37610 2544
rect 37554 2488 37556 2508
rect 37556 2488 37608 2508
rect 37608 2488 37610 2508
rect 38290 6704 38346 6760
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 24117 36954 24183 36957
rect 20118 36952 24183 36954
rect 20118 36896 24122 36952
rect 24178 36896 24183 36952
rect 20118 36894 24183 36896
rect 17677 36818 17743 36821
rect 20118 36818 20178 36894
rect 24117 36891 24183 36894
rect 24669 36954 24735 36957
rect 28165 36954 28231 36957
rect 24669 36952 28231 36954
rect 24669 36896 24674 36952
rect 24730 36896 28170 36952
rect 28226 36896 28231 36952
rect 24669 36894 28231 36896
rect 24669 36891 24735 36894
rect 28165 36891 28231 36894
rect 17677 36816 20178 36818
rect 17677 36760 17682 36816
rect 17738 36760 20178 36816
rect 17677 36758 20178 36760
rect 23381 36818 23447 36821
rect 25773 36818 25839 36821
rect 26325 36818 26391 36821
rect 23381 36816 26391 36818
rect 23381 36760 23386 36816
rect 23442 36760 25778 36816
rect 25834 36760 26330 36816
rect 26386 36760 26391 36816
rect 23381 36758 26391 36760
rect 17677 36755 17743 36758
rect 23381 36755 23447 36758
rect 25773 36755 25839 36758
rect 26325 36755 26391 36758
rect 23381 36682 23447 36685
rect 25405 36682 25471 36685
rect 23381 36680 25471 36682
rect 23381 36624 23386 36680
rect 23442 36624 25410 36680
rect 25466 36624 25471 36680
rect 23381 36622 25471 36624
rect 23381 36619 23447 36622
rect 25405 36619 25471 36622
rect 21030 36484 21036 36548
rect 21100 36546 21106 36548
rect 21173 36546 21239 36549
rect 21100 36544 21239 36546
rect 21100 36488 21178 36544
rect 21234 36488 21239 36544
rect 21100 36486 21239 36488
rect 21100 36484 21106 36486
rect 21173 36483 21239 36486
rect 22369 36546 22435 36549
rect 26141 36546 26207 36549
rect 22369 36544 26207 36546
rect 22369 36488 22374 36544
rect 22430 36488 26146 36544
rect 26202 36488 26207 36544
rect 22369 36486 26207 36488
rect 22369 36483 22435 36486
rect 26141 36483 26207 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 21081 36410 21147 36413
rect 33961 36410 34027 36413
rect 21081 36408 34027 36410
rect 21081 36352 21086 36408
rect 21142 36352 33966 36408
rect 34022 36352 34027 36408
rect 21081 36350 34027 36352
rect 21081 36347 21147 36350
rect 33961 36347 34027 36350
rect 21725 36274 21791 36277
rect 26969 36274 27035 36277
rect 21725 36272 27035 36274
rect 21725 36216 21730 36272
rect 21786 36216 26974 36272
rect 27030 36216 27035 36272
rect 21725 36214 27035 36216
rect 21725 36211 21791 36214
rect 26969 36211 27035 36214
rect 10225 36138 10291 36141
rect 19057 36138 19123 36141
rect 24577 36138 24643 36141
rect 30281 36138 30347 36141
rect 10225 36136 20178 36138
rect 10225 36080 10230 36136
rect 10286 36080 19062 36136
rect 19118 36080 20178 36136
rect 10225 36078 20178 36080
rect 10225 36075 10291 36078
rect 19057 36075 19123 36078
rect 20118 36002 20178 36078
rect 24577 36136 30347 36138
rect 24577 36080 24582 36136
rect 24638 36080 30286 36136
rect 30342 36080 30347 36136
rect 24577 36078 30347 36080
rect 24577 36075 24643 36078
rect 30281 36075 30347 36078
rect 24301 36002 24367 36005
rect 36537 36004 36603 36005
rect 20118 36000 24367 36002
rect 20118 35944 24306 36000
rect 24362 35944 24367 36000
rect 20118 35942 24367 35944
rect 24301 35939 24367 35942
rect 36486 35940 36492 36004
rect 36556 36002 36603 36004
rect 36556 36000 36648 36002
rect 36598 35944 36648 36000
rect 36556 35942 36648 35944
rect 36556 35940 36603 35942
rect 36537 35939 36603 35940
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 22737 35866 22803 35869
rect 25129 35866 25195 35869
rect 26233 35866 26299 35869
rect 22737 35864 26299 35866
rect 22737 35808 22742 35864
rect 22798 35808 25134 35864
rect 25190 35808 26238 35864
rect 26294 35808 26299 35864
rect 22737 35806 26299 35808
rect 22737 35803 22803 35806
rect 25129 35803 25195 35806
rect 26233 35803 26299 35806
rect 19333 35730 19399 35733
rect 34605 35730 34671 35733
rect 19333 35728 34671 35730
rect 19333 35672 19338 35728
rect 19394 35672 34610 35728
rect 34666 35672 34671 35728
rect 19333 35670 34671 35672
rect 19333 35667 19399 35670
rect 34605 35667 34671 35670
rect 23381 35458 23447 35461
rect 25405 35458 25471 35461
rect 23381 35456 25471 35458
rect 23381 35400 23386 35456
rect 23442 35400 25410 35456
rect 25466 35400 25471 35456
rect 23381 35398 25471 35400
rect 23381 35395 23447 35398
rect 25405 35395 25471 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 12433 35322 12499 35325
rect 28993 35322 29059 35325
rect 12433 35320 29059 35322
rect 12433 35264 12438 35320
rect 12494 35264 28998 35320
rect 29054 35264 29059 35320
rect 12433 35262 29059 35264
rect 12433 35259 12499 35262
rect 28993 35259 29059 35262
rect 21633 35186 21699 35189
rect 31385 35186 31451 35189
rect 21633 35184 31451 35186
rect 21633 35128 21638 35184
rect 21694 35128 31390 35184
rect 31446 35128 31451 35184
rect 21633 35126 31451 35128
rect 21633 35123 21699 35126
rect 31385 35123 31451 35126
rect 19977 35050 20043 35053
rect 34513 35050 34579 35053
rect 19977 35048 34579 35050
rect 19977 34992 19982 35048
rect 20038 34992 34518 35048
rect 34574 34992 34579 35048
rect 19977 34990 34579 34992
rect 19977 34987 20043 34990
rect 34513 34987 34579 34990
rect 34605 34916 34671 34917
rect 34605 34914 34652 34916
rect 34560 34912 34652 34914
rect 34560 34856 34610 34912
rect 34560 34854 34652 34856
rect 34605 34852 34652 34854
rect 34716 34852 34722 34916
rect 34605 34851 34671 34852
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 23381 34778 23447 34781
rect 31845 34778 31911 34781
rect 23381 34776 31911 34778
rect 23381 34720 23386 34776
rect 23442 34720 31850 34776
rect 31906 34720 31911 34776
rect 23381 34718 31911 34720
rect 23381 34715 23447 34718
rect 31845 34715 31911 34718
rect 12065 34642 12131 34645
rect 26969 34642 27035 34645
rect 12065 34640 27035 34642
rect 12065 34584 12070 34640
rect 12126 34584 26974 34640
rect 27030 34584 27035 34640
rect 12065 34582 27035 34584
rect 12065 34579 12131 34582
rect 26969 34579 27035 34582
rect 24117 34506 24183 34509
rect 36261 34506 36327 34509
rect 24117 34504 36327 34506
rect 24117 34448 24122 34504
rect 24178 34448 36266 34504
rect 36322 34448 36327 34504
rect 24117 34446 36327 34448
rect 24117 34443 24183 34446
rect 36261 34443 36327 34446
rect 22185 34370 22251 34373
rect 29177 34370 29243 34373
rect 22185 34368 29243 34370
rect 22185 34312 22190 34368
rect 22246 34312 29182 34368
rect 29238 34312 29243 34368
rect 22185 34310 29243 34312
rect 22185 34307 22251 34310
rect 29177 34307 29243 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 12249 34234 12315 34237
rect 27797 34234 27863 34237
rect 12249 34232 27863 34234
rect 12249 34176 12254 34232
rect 12310 34176 27802 34232
rect 27858 34176 27863 34232
rect 12249 34174 27863 34176
rect 12249 34171 12315 34174
rect 27797 34171 27863 34174
rect 24577 34098 24643 34101
rect 31661 34098 31727 34101
rect 24577 34096 31727 34098
rect 24577 34040 24582 34096
rect 24638 34040 31666 34096
rect 31722 34040 31727 34096
rect 24577 34038 31727 34040
rect 24577 34035 24643 34038
rect 31661 34035 31727 34038
rect 18321 33962 18387 33965
rect 34513 33962 34579 33965
rect 18321 33960 34579 33962
rect 18321 33904 18326 33960
rect 18382 33904 34518 33960
rect 34574 33904 34579 33960
rect 18321 33902 34579 33904
rect 18321 33899 18387 33902
rect 34513 33899 34579 33902
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 22737 33554 22803 33557
rect 33041 33554 33107 33557
rect 22737 33552 33107 33554
rect 22737 33496 22742 33552
rect 22798 33496 33046 33552
rect 33102 33496 33107 33552
rect 22737 33494 33107 33496
rect 22737 33491 22803 33494
rect 33041 33491 33107 33494
rect 24117 33282 24183 33285
rect 26325 33282 26391 33285
rect 24117 33280 26391 33282
rect 24117 33224 24122 33280
rect 24178 33224 26330 33280
rect 26386 33224 26391 33280
rect 24117 33222 26391 33224
rect 24117 33219 24183 33222
rect 26325 33219 26391 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 20805 33146 20871 33149
rect 28993 33146 29059 33149
rect 20805 33144 29059 33146
rect 20805 33088 20810 33144
rect 20866 33088 28998 33144
rect 29054 33088 29059 33144
rect 20805 33086 29059 33088
rect 20805 33083 20871 33086
rect 28993 33083 29059 33086
rect 22737 33010 22803 33013
rect 23238 33010 23244 33012
rect 22737 33008 23244 33010
rect 22737 32952 22742 33008
rect 22798 32952 23244 33008
rect 22737 32950 23244 32952
rect 22737 32947 22803 32950
rect 23238 32948 23244 32950
rect 23308 32948 23314 33012
rect 22737 32874 22803 32877
rect 33317 32874 33383 32877
rect 22737 32872 33383 32874
rect 22737 32816 22742 32872
rect 22798 32816 33322 32872
rect 33378 32816 33383 32872
rect 22737 32814 33383 32816
rect 22737 32811 22803 32814
rect 33317 32811 33383 32814
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 23381 32602 23447 32605
rect 27245 32602 27311 32605
rect 23381 32600 27311 32602
rect 23381 32544 23386 32600
rect 23442 32544 27250 32600
rect 27306 32544 27311 32600
rect 23381 32542 27311 32544
rect 23381 32539 23447 32542
rect 27245 32539 27311 32542
rect 13261 32330 13327 32333
rect 14825 32330 14891 32333
rect 31017 32330 31083 32333
rect 13261 32328 31083 32330
rect 13261 32272 13266 32328
rect 13322 32272 14830 32328
rect 14886 32272 31022 32328
rect 31078 32272 31083 32328
rect 13261 32270 31083 32272
rect 13261 32267 13327 32270
rect 14825 32267 14891 32270
rect 31017 32267 31083 32270
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 13629 31786 13695 31789
rect 24393 31786 24459 31789
rect 13629 31784 24459 31786
rect 13629 31728 13634 31784
rect 13690 31728 24398 31784
rect 24454 31728 24459 31784
rect 13629 31726 24459 31728
rect 13629 31723 13695 31726
rect 24393 31723 24459 31726
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 16849 31106 16915 31109
rect 17677 31106 17743 31109
rect 28349 31106 28415 31109
rect 16849 31104 28415 31106
rect 16849 31048 16854 31104
rect 16910 31048 17682 31104
rect 17738 31048 28354 31104
rect 28410 31048 28415 31104
rect 16849 31046 28415 31048
rect 16849 31043 16915 31046
rect 17677 31043 17743 31046
rect 28349 31043 28415 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 16481 30290 16547 30293
rect 19057 30290 19123 30293
rect 16481 30288 19123 30290
rect 16481 30232 16486 30288
rect 16542 30232 19062 30288
rect 19118 30232 19123 30288
rect 16481 30230 19123 30232
rect 16481 30227 16547 30230
rect 19057 30227 19123 30230
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 13537 29746 13603 29749
rect 24669 29746 24735 29749
rect 13537 29744 24735 29746
rect 13537 29688 13542 29744
rect 13598 29688 24674 29744
rect 24730 29688 24735 29744
rect 13537 29686 24735 29688
rect 13537 29683 13603 29686
rect 24669 29683 24735 29686
rect 14273 29610 14339 29613
rect 29545 29610 29611 29613
rect 14273 29608 29611 29610
rect 14273 29552 14278 29608
rect 14334 29552 29550 29608
rect 29606 29552 29611 29608
rect 14273 29550 29611 29552
rect 14273 29547 14339 29550
rect 29545 29547 29611 29550
rect 20989 29474 21055 29477
rect 24393 29474 24459 29477
rect 20989 29472 24459 29474
rect 20989 29416 20994 29472
rect 21050 29416 24398 29472
rect 24454 29416 24459 29472
rect 20989 29414 24459 29416
rect 20989 29411 21055 29414
rect 24393 29411 24459 29414
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 20529 29338 20595 29341
rect 21817 29338 21883 29341
rect 20529 29336 21883 29338
rect 20529 29280 20534 29336
rect 20590 29280 21822 29336
rect 21878 29280 21883 29336
rect 20529 29278 21883 29280
rect 20529 29275 20595 29278
rect 21817 29275 21883 29278
rect 13169 29202 13235 29205
rect 25037 29202 25103 29205
rect 13169 29200 25103 29202
rect 13169 29144 13174 29200
rect 13230 29144 25042 29200
rect 25098 29144 25103 29200
rect 13169 29142 25103 29144
rect 13169 29139 13235 29142
rect 25037 29139 25103 29142
rect 12341 29066 12407 29069
rect 27613 29066 27679 29069
rect 12341 29064 27679 29066
rect 12341 29008 12346 29064
rect 12402 29008 27618 29064
rect 27674 29008 27679 29064
rect 12341 29006 27679 29008
rect 12341 29003 12407 29006
rect 27613 29003 27679 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 12341 28522 12407 28525
rect 26969 28522 27035 28525
rect 12341 28520 27035 28522
rect 12341 28464 12346 28520
rect 12402 28464 26974 28520
rect 27030 28464 27035 28520
rect 12341 28462 27035 28464
rect 12341 28459 12407 28462
rect 26969 28459 27035 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 9949 28114 10015 28117
rect 24853 28114 24919 28117
rect 9949 28112 24919 28114
rect 9949 28056 9954 28112
rect 10010 28056 24858 28112
rect 24914 28056 24919 28112
rect 9949 28054 24919 28056
rect 9949 28051 10015 28054
rect 24853 28051 24919 28054
rect 16849 27978 16915 27981
rect 34605 27978 34671 27981
rect 16849 27976 34671 27978
rect 16849 27920 16854 27976
rect 16910 27920 34610 27976
rect 34666 27920 34671 27976
rect 16849 27918 34671 27920
rect 16849 27915 16915 27918
rect 34605 27915 34671 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 18689 27570 18755 27573
rect 31753 27570 31819 27573
rect 18689 27568 31819 27570
rect 18689 27512 18694 27568
rect 18750 27512 31758 27568
rect 31814 27512 31819 27568
rect 18689 27510 31819 27512
rect 18689 27507 18755 27510
rect 31753 27507 31819 27510
rect 9489 27434 9555 27437
rect 24853 27434 24919 27437
rect 9489 27432 24919 27434
rect 9489 27376 9494 27432
rect 9550 27376 24858 27432
rect 24914 27376 24919 27432
rect 9489 27374 24919 27376
rect 9489 27371 9555 27374
rect 24853 27371 24919 27374
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 16389 27026 16455 27029
rect 21449 27026 21515 27029
rect 16389 27024 21515 27026
rect 16389 26968 16394 27024
rect 16450 26968 21454 27024
rect 21510 26968 21515 27024
rect 16389 26966 21515 26968
rect 16389 26963 16455 26966
rect 21449 26963 21515 26966
rect 10225 26890 10291 26893
rect 25221 26890 25287 26893
rect 10225 26888 25287 26890
rect 10225 26832 10230 26888
rect 10286 26832 25226 26888
rect 25282 26832 25287 26888
rect 10225 26830 25287 26832
rect 10225 26827 10291 26830
rect 25221 26827 25287 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19517 26482 19583 26485
rect 20621 26482 20687 26485
rect 19517 26480 20687 26482
rect 19517 26424 19522 26480
rect 19578 26424 20626 26480
rect 20682 26424 20687 26480
rect 19517 26422 20687 26424
rect 19517 26419 19583 26422
rect 20621 26419 20687 26422
rect 11881 26346 11947 26349
rect 27613 26346 27679 26349
rect 11881 26344 27679 26346
rect 11881 26288 11886 26344
rect 11942 26288 27618 26344
rect 27674 26288 27679 26344
rect 11881 26286 27679 26288
rect 11881 26283 11947 26286
rect 27613 26283 27679 26286
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 31201 26074 31267 26077
rect 22050 26072 31267 26074
rect 22050 26016 31206 26072
rect 31262 26016 31267 26072
rect 22050 26014 31267 26016
rect 17033 25938 17099 25941
rect 22050 25938 22110 26014
rect 31201 26011 31267 26014
rect 17033 25936 22110 25938
rect 17033 25880 17038 25936
rect 17094 25880 22110 25936
rect 17033 25878 22110 25880
rect 22553 25938 22619 25941
rect 28901 25938 28967 25941
rect 22553 25936 28967 25938
rect 22553 25880 22558 25936
rect 22614 25880 28906 25936
rect 28962 25880 28967 25936
rect 22553 25878 28967 25880
rect 17033 25875 17099 25878
rect 22553 25875 22619 25878
rect 28901 25875 28967 25878
rect 36077 25802 36143 25805
rect 22050 25800 36143 25802
rect 22050 25744 36082 25800
rect 36138 25744 36143 25800
rect 22050 25742 36143 25744
rect 16665 25666 16731 25669
rect 22050 25666 22110 25742
rect 36077 25739 36143 25742
rect 16665 25664 22110 25666
rect 16665 25608 16670 25664
rect 16726 25608 22110 25664
rect 16665 25606 22110 25608
rect 16665 25603 16731 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 18413 25530 18479 25533
rect 27981 25530 28047 25533
rect 18413 25528 28047 25530
rect 18413 25472 18418 25528
rect 18474 25472 27986 25528
rect 28042 25472 28047 25528
rect 18413 25470 28047 25472
rect 18413 25467 18479 25470
rect 27981 25467 28047 25470
rect 10225 25394 10291 25397
rect 24393 25394 24459 25397
rect 10225 25392 24459 25394
rect 10225 25336 10230 25392
rect 10286 25336 24398 25392
rect 24454 25336 24459 25392
rect 10225 25334 24459 25336
rect 10225 25331 10291 25334
rect 24393 25331 24459 25334
rect 8845 25258 8911 25261
rect 23657 25258 23723 25261
rect 8845 25256 23723 25258
rect 8845 25200 8850 25256
rect 8906 25200 23662 25256
rect 23718 25200 23723 25256
rect 8845 25198 23723 25200
rect 8845 25195 8911 25198
rect 23657 25195 23723 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 20437 24850 20503 24853
rect 27705 24850 27771 24853
rect 20437 24848 27771 24850
rect 20437 24792 20442 24848
rect 20498 24792 27710 24848
rect 27766 24792 27771 24848
rect 20437 24790 27771 24792
rect 20437 24787 20503 24790
rect 27705 24787 27771 24790
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 20069 23762 20135 23765
rect 30925 23762 30991 23765
rect 20069 23760 30991 23762
rect 20069 23704 20074 23760
rect 20130 23704 30930 23760
rect 30986 23704 30991 23760
rect 20069 23702 30991 23704
rect 20069 23699 20135 23702
rect 30925 23699 30991 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 32305 22810 32371 22813
rect 36905 22810 36971 22813
rect 32305 22808 36971 22810
rect 32305 22752 32310 22808
rect 32366 22752 36910 22808
rect 36966 22752 36971 22808
rect 32305 22750 36971 22752
rect 32305 22747 32371 22750
rect 36905 22747 36971 22750
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 36445 19956 36511 19957
rect 36445 19954 36492 19956
rect 36400 19952 36492 19954
rect 36400 19896 36450 19952
rect 36400 19894 36492 19896
rect 36445 19892 36492 19894
rect 36556 19892 36562 19956
rect 36445 19891 36511 19892
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 18321 17234 18387 17237
rect 19374 17234 19380 17236
rect 18321 17232 19380 17234
rect 18321 17176 18326 17232
rect 18382 17176 19380 17232
rect 18321 17174 19380 17176
rect 18321 17171 18387 17174
rect 19374 17172 19380 17174
rect 19444 17172 19450 17236
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 23238 15132 23244 15196
rect 23308 15194 23314 15196
rect 24945 15194 25011 15197
rect 23308 15192 25011 15194
rect 23308 15136 24950 15192
rect 25006 15136 25011 15192
rect 23308 15134 25011 15136
rect 23308 15132 23314 15134
rect 24945 15131 25011 15134
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 20621 14650 20687 14653
rect 21030 14650 21036 14652
rect 20621 14648 21036 14650
rect 20621 14592 20626 14648
rect 20682 14592 21036 14648
rect 20621 14590 21036 14592
rect 20621 14587 20687 14590
rect 21030 14588 21036 14590
rect 21100 14588 21106 14652
rect 26417 14650 26483 14653
rect 34646 14650 34652 14652
rect 26417 14648 34652 14650
rect 26417 14592 26422 14648
rect 26478 14592 34652 14648
rect 26417 14590 34652 14592
rect 26417 14587 26483 14590
rect 34646 14588 34652 14590
rect 34716 14588 34722 14652
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 18689 13836 18755 13837
rect 18638 13834 18644 13836
rect 18598 13774 18644 13834
rect 18708 13832 18755 13836
rect 18750 13776 18755 13832
rect 18638 13772 18644 13774
rect 18708 13772 18755 13776
rect 18689 13771 18755 13772
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 16205 13426 16271 13429
rect 24485 13426 24551 13429
rect 16205 13424 24551 13426
rect 16205 13368 16210 13424
rect 16266 13368 24490 13424
rect 24546 13368 24551 13424
rect 16205 13366 24551 13368
rect 16205 13363 16271 13366
rect 24485 13363 24551 13366
rect 20069 13290 20135 13293
rect 29545 13290 29611 13293
rect 20069 13288 29611 13290
rect 20069 13232 20074 13288
rect 20130 13232 29550 13288
rect 29606 13232 29611 13288
rect 20069 13230 29611 13232
rect 20069 13227 20135 13230
rect 29545 13227 29611 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 15285 12338 15351 12341
rect 21633 12338 21699 12341
rect 15285 12336 21699 12338
rect 15285 12280 15290 12336
rect 15346 12280 21638 12336
rect 21694 12280 21699 12336
rect 15285 12278 21699 12280
rect 15285 12275 15351 12278
rect 21633 12275 21699 12278
rect 20621 12202 20687 12205
rect 27705 12202 27771 12205
rect 20621 12200 27771 12202
rect 20621 12144 20626 12200
rect 20682 12144 27710 12200
rect 27766 12144 27771 12200
rect 20621 12142 27771 12144
rect 20621 12139 20687 12142
rect 27705 12139 27771 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 16481 11658 16547 11661
rect 23381 11658 23447 11661
rect 16481 11656 23447 11658
rect 16481 11600 16486 11656
rect 16542 11600 23386 11656
rect 23442 11600 23447 11656
rect 16481 11598 23447 11600
rect 16481 11595 16547 11598
rect 23381 11595 23447 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 15193 11250 15259 11253
rect 17953 11250 18019 11253
rect 15193 11248 18019 11250
rect 15193 11192 15198 11248
rect 15254 11192 17958 11248
rect 18014 11192 18019 11248
rect 15193 11190 18019 11192
rect 15193 11187 15259 11190
rect 17953 11187 18019 11190
rect 16665 11114 16731 11117
rect 17033 11114 17099 11117
rect 21725 11114 21791 11117
rect 16665 11112 21791 11114
rect 16665 11056 16670 11112
rect 16726 11056 17038 11112
rect 17094 11056 21730 11112
rect 21786 11056 21791 11112
rect 16665 11054 21791 11056
rect 16665 11051 16731 11054
rect 17033 11051 17099 11054
rect 21725 11051 21791 11054
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 11697 10570 11763 10573
rect 26233 10570 26299 10573
rect 11697 10568 26299 10570
rect 11697 10512 11702 10568
rect 11758 10512 26238 10568
rect 26294 10512 26299 10568
rect 11697 10510 26299 10512
rect 11697 10507 11763 10510
rect 26233 10507 26299 10510
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 10869 10162 10935 10165
rect 23381 10162 23447 10165
rect 10869 10160 23447 10162
rect 10869 10104 10874 10160
rect 10930 10104 23386 10160
rect 23442 10104 23447 10160
rect 10869 10102 23447 10104
rect 10869 10099 10935 10102
rect 23381 10099 23447 10102
rect 14825 10026 14891 10029
rect 16297 10026 16363 10029
rect 21817 10026 21883 10029
rect 14825 10024 21883 10026
rect 14825 9968 14830 10024
rect 14886 9968 16302 10024
rect 16358 9968 21822 10024
rect 21878 9968 21883 10024
rect 14825 9966 21883 9968
rect 14825 9963 14891 9966
rect 16297 9963 16363 9966
rect 21817 9963 21883 9966
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 12801 9482 12867 9485
rect 25221 9482 25287 9485
rect 12801 9480 25287 9482
rect 12801 9424 12806 9480
rect 12862 9424 25226 9480
rect 25282 9424 25287 9480
rect 12801 9422 25287 9424
rect 12801 9419 12867 9422
rect 25221 9419 25287 9422
rect 24945 9346 25011 9349
rect 29361 9346 29427 9349
rect 24945 9344 29427 9346
rect 24945 9288 24950 9344
rect 25006 9288 29366 9344
rect 29422 9288 29427 9344
rect 24945 9286 29427 9288
rect 24945 9283 25011 9286
rect 29361 9283 29427 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 16941 9210 17007 9213
rect 26417 9210 26483 9213
rect 16941 9208 26483 9210
rect 16941 9152 16946 9208
rect 17002 9152 26422 9208
rect 26478 9152 26483 9208
rect 16941 9150 26483 9152
rect 16941 9147 17007 9150
rect 26417 9147 26483 9150
rect 13721 9074 13787 9077
rect 21081 9074 21147 9077
rect 13721 9072 21147 9074
rect 13721 9016 13726 9072
rect 13782 9016 21086 9072
rect 21142 9016 21147 9072
rect 13721 9014 21147 9016
rect 13721 9011 13787 9014
rect 21081 9011 21147 9014
rect 10225 8938 10291 8941
rect 24025 8938 24091 8941
rect 10225 8936 24091 8938
rect 10225 8880 10230 8936
rect 10286 8880 24030 8936
rect 24086 8880 24091 8936
rect 10225 8878 24091 8880
rect 10225 8875 10291 8878
rect 24025 8875 24091 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 20437 8530 20503 8533
rect 26233 8530 26299 8533
rect 20437 8528 26299 8530
rect 20437 8472 20442 8528
rect 20498 8472 26238 8528
rect 26294 8472 26299 8528
rect 20437 8470 26299 8472
rect 20437 8467 20503 8470
rect 26233 8467 26299 8470
rect 20253 8394 20319 8397
rect 37365 8394 37431 8397
rect 20253 8392 37431 8394
rect 20253 8336 20258 8392
rect 20314 8336 37370 8392
rect 37426 8336 37431 8392
rect 20253 8334 37431 8336
rect 20253 8331 20319 8334
rect 37365 8331 37431 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 15101 7850 15167 7853
rect 22001 7850 22067 7853
rect 15101 7848 22067 7850
rect 15101 7792 15106 7848
rect 15162 7792 22006 7848
rect 22062 7792 22067 7848
rect 15101 7790 22067 7792
rect 15101 7787 15167 7790
rect 22001 7787 22067 7790
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 17401 7442 17467 7445
rect 30373 7442 30439 7445
rect 17401 7440 30439 7442
rect 17401 7384 17406 7440
rect 17462 7384 30378 7440
rect 30434 7384 30439 7440
rect 17401 7382 30439 7384
rect 17401 7379 17467 7382
rect 30373 7379 30439 7382
rect 17953 7306 18019 7309
rect 22277 7306 22343 7309
rect 17953 7304 22343 7306
rect 17953 7248 17958 7304
rect 18014 7248 22282 7304
rect 22338 7248 22343 7304
rect 17953 7246 22343 7248
rect 17953 7243 18019 7246
rect 22277 7243 22343 7246
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 11697 7034 11763 7037
rect 23565 7034 23631 7037
rect 11697 7032 23631 7034
rect 11697 6976 11702 7032
rect 11758 6976 23570 7032
rect 23626 6976 23631 7032
rect 11697 6974 23631 6976
rect 11697 6971 11763 6974
rect 23565 6971 23631 6974
rect 19374 6836 19380 6900
rect 19444 6898 19450 6900
rect 22369 6898 22435 6901
rect 19444 6896 22435 6898
rect 19444 6840 22374 6896
rect 22430 6840 22435 6896
rect 19444 6838 22435 6840
rect 19444 6836 19450 6838
rect 22369 6835 22435 6838
rect 13353 6762 13419 6765
rect 21633 6762 21699 6765
rect 13353 6760 21699 6762
rect 13353 6704 13358 6760
rect 13414 6704 21638 6760
rect 21694 6704 21699 6760
rect 13353 6702 21699 6704
rect 13353 6699 13419 6702
rect 21633 6699 21699 6702
rect 37549 6762 37615 6765
rect 38285 6762 38351 6765
rect 37549 6760 38351 6762
rect 37549 6704 37554 6760
rect 37610 6704 38290 6760
rect 38346 6704 38351 6760
rect 37549 6702 38351 6704
rect 37549 6699 37615 6702
rect 38285 6699 38351 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 19057 6354 19123 6357
rect 28993 6354 29059 6357
rect 19057 6352 29059 6354
rect 19057 6296 19062 6352
rect 19118 6296 28998 6352
rect 29054 6296 29059 6352
rect 19057 6294 29059 6296
rect 19057 6291 19123 6294
rect 28993 6291 29059 6294
rect 15745 6218 15811 6221
rect 37457 6218 37523 6221
rect 15745 6216 37523 6218
rect 15745 6160 15750 6216
rect 15806 6160 37462 6216
rect 37518 6160 37523 6216
rect 15745 6158 37523 6160
rect 15745 6155 15811 6158
rect 37457 6155 37523 6158
rect 18689 6082 18755 6085
rect 26141 6082 26207 6085
rect 18689 6080 26207 6082
rect 18689 6024 18694 6080
rect 18750 6024 26146 6080
rect 26202 6024 26207 6080
rect 18689 6022 26207 6024
rect 18689 6019 18755 6022
rect 26141 6019 26207 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 12893 5946 12959 5949
rect 22645 5946 22711 5949
rect 12893 5944 22711 5946
rect 12893 5888 12898 5944
rect 12954 5888 22650 5944
rect 22706 5888 22711 5944
rect 12893 5886 22711 5888
rect 12893 5883 12959 5886
rect 22645 5883 22711 5886
rect 11053 5810 11119 5813
rect 16941 5810 17007 5813
rect 11053 5808 17007 5810
rect 11053 5752 11058 5808
rect 11114 5752 16946 5808
rect 17002 5752 17007 5808
rect 11053 5750 17007 5752
rect 11053 5747 11119 5750
rect 16941 5747 17007 5750
rect 17585 5810 17651 5813
rect 27613 5810 27679 5813
rect 17585 5808 27679 5810
rect 17585 5752 17590 5808
rect 17646 5752 27618 5808
rect 27674 5752 27679 5808
rect 17585 5750 27679 5752
rect 17585 5747 17651 5750
rect 27613 5747 27679 5750
rect 9673 5674 9739 5677
rect 20805 5674 20871 5677
rect 9673 5672 20871 5674
rect 9673 5616 9678 5672
rect 9734 5616 20810 5672
rect 20866 5616 20871 5672
rect 9673 5614 20871 5616
rect 9673 5611 9739 5614
rect 20805 5611 20871 5614
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 10501 5266 10567 5269
rect 21817 5266 21883 5269
rect 10501 5264 21883 5266
rect 10501 5208 10506 5264
rect 10562 5208 21822 5264
rect 21878 5208 21883 5264
rect 10501 5206 21883 5208
rect 10501 5203 10567 5206
rect 21817 5203 21883 5206
rect 15837 5130 15903 5133
rect 26417 5130 26483 5133
rect 15837 5128 26483 5130
rect 15837 5072 15842 5128
rect 15898 5072 26422 5128
rect 26478 5072 26483 5128
rect 15837 5070 26483 5072
rect 15837 5067 15903 5070
rect 26417 5067 26483 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 13721 4586 13787 4589
rect 22369 4586 22435 4589
rect 13721 4584 22435 4586
rect 13721 4528 13726 4584
rect 13782 4528 22374 4584
rect 22430 4528 22435 4584
rect 13721 4526 22435 4528
rect 13721 4523 13787 4526
rect 22369 4523 22435 4526
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 18137 4314 18203 4317
rect 20529 4314 20595 4317
rect 28441 4314 28507 4317
rect 18137 4312 19442 4314
rect 18137 4256 18142 4312
rect 18198 4256 19442 4312
rect 18137 4254 19442 4256
rect 18137 4251 18203 4254
rect 12249 4178 12315 4181
rect 15377 4178 15443 4181
rect 12249 4176 15443 4178
rect 12249 4120 12254 4176
rect 12310 4120 15382 4176
rect 15438 4120 15443 4176
rect 12249 4118 15443 4120
rect 12249 4115 12315 4118
rect 15377 4115 15443 4118
rect 18229 4178 18295 4181
rect 19190 4178 19196 4180
rect 18229 4176 19196 4178
rect 18229 4120 18234 4176
rect 18290 4120 19196 4176
rect 18229 4118 19196 4120
rect 18229 4115 18295 4118
rect 19190 4116 19196 4118
rect 19260 4116 19266 4180
rect 19382 4178 19442 4254
rect 20529 4312 28507 4314
rect 20529 4256 20534 4312
rect 20590 4256 28446 4312
rect 28502 4256 28507 4312
rect 20529 4254 28507 4256
rect 20529 4251 20595 4254
rect 28441 4251 28507 4254
rect 24577 4178 24643 4181
rect 19382 4176 24643 4178
rect 19382 4120 24582 4176
rect 24638 4120 24643 4176
rect 19382 4118 24643 4120
rect 24577 4115 24643 4118
rect 10593 4042 10659 4045
rect 12709 4042 12775 4045
rect 10593 4040 12775 4042
rect 10593 3984 10598 4040
rect 10654 3984 12714 4040
rect 12770 3984 12775 4040
rect 10593 3982 12775 3984
rect 10593 3979 10659 3982
rect 12709 3979 12775 3982
rect 13169 4042 13235 4045
rect 13537 4042 13603 4045
rect 20805 4042 20871 4045
rect 13169 4040 20871 4042
rect 13169 3984 13174 4040
rect 13230 3984 13542 4040
rect 13598 3984 20810 4040
rect 20866 3984 20871 4040
rect 13169 3982 20871 3984
rect 13169 3979 13235 3982
rect 13537 3979 13603 3982
rect 20805 3979 20871 3982
rect 9397 3906 9463 3909
rect 13721 3906 13787 3909
rect 21633 3906 21699 3909
rect 9397 3904 13787 3906
rect 9397 3848 9402 3904
rect 9458 3848 13726 3904
rect 13782 3848 13787 3904
rect 9397 3846 13787 3848
rect 9397 3843 9463 3846
rect 13721 3843 13787 3846
rect 16990 3904 21699 3906
rect 16990 3848 21638 3904
rect 21694 3848 21699 3904
rect 16990 3846 21699 3848
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 7189 3770 7255 3773
rect 10409 3770 10475 3773
rect 12341 3770 12407 3773
rect 16990 3770 17050 3846
rect 21633 3843 21699 3846
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 7189 3768 17050 3770
rect 7189 3712 7194 3768
rect 7250 3712 10414 3768
rect 10470 3712 12346 3768
rect 12402 3712 17050 3768
rect 7189 3710 17050 3712
rect 19241 3770 19307 3773
rect 28073 3770 28139 3773
rect 19241 3768 28139 3770
rect 19241 3712 19246 3768
rect 19302 3712 28078 3768
rect 28134 3712 28139 3768
rect 19241 3710 28139 3712
rect 7189 3707 7255 3710
rect 10409 3707 10475 3710
rect 12341 3707 12407 3710
rect 19241 3707 19307 3710
rect 28073 3707 28139 3710
rect 28993 3770 29059 3773
rect 31753 3770 31819 3773
rect 28993 3768 31819 3770
rect 28993 3712 28998 3768
rect 29054 3712 31758 3768
rect 31814 3712 31819 3768
rect 28993 3710 31819 3712
rect 28993 3707 29059 3710
rect 31753 3707 31819 3710
rect 6177 3634 6243 3637
rect 9121 3634 9187 3637
rect 11973 3634 12039 3637
rect 13537 3634 13603 3637
rect 6177 3632 9322 3634
rect 6177 3576 6182 3632
rect 6238 3576 9126 3632
rect 9182 3576 9322 3632
rect 6177 3574 9322 3576
rect 6177 3571 6243 3574
rect 9121 3571 9187 3574
rect 9262 3498 9322 3574
rect 11973 3632 13603 3634
rect 11973 3576 11978 3632
rect 12034 3576 13542 3632
rect 13598 3576 13603 3632
rect 11973 3574 13603 3576
rect 11973 3571 12039 3574
rect 13537 3571 13603 3574
rect 19374 3572 19380 3636
rect 19444 3634 19450 3636
rect 19701 3634 19767 3637
rect 20437 3634 20503 3637
rect 19444 3632 20503 3634
rect 19444 3576 19706 3632
rect 19762 3576 20442 3632
rect 20498 3576 20503 3632
rect 19444 3574 20503 3576
rect 19444 3572 19450 3574
rect 19701 3571 19767 3574
rect 20437 3571 20503 3574
rect 20805 3634 20871 3637
rect 25865 3634 25931 3637
rect 20805 3632 25931 3634
rect 20805 3576 20810 3632
rect 20866 3576 25870 3632
rect 25926 3576 25931 3632
rect 20805 3574 25931 3576
rect 20805 3571 20871 3574
rect 25865 3571 25931 3574
rect 25497 3498 25563 3501
rect 9262 3496 25563 3498
rect 9262 3440 25502 3496
rect 25558 3440 25563 3496
rect 9262 3438 25563 3440
rect 25497 3435 25563 3438
rect 35985 3498 36051 3501
rect 36997 3498 37063 3501
rect 35985 3496 37063 3498
rect 35985 3440 35990 3496
rect 36046 3440 37002 3496
rect 37058 3440 37063 3496
rect 35985 3438 37063 3440
rect 35985 3435 36051 3438
rect 36997 3435 37063 3438
rect 11513 3362 11579 3365
rect 12157 3362 12223 3365
rect 11513 3360 12223 3362
rect 11513 3304 11518 3360
rect 11574 3304 12162 3360
rect 12218 3304 12223 3360
rect 11513 3302 12223 3304
rect 11513 3299 11579 3302
rect 12157 3299 12223 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 9949 3226 10015 3229
rect 16297 3226 16363 3229
rect 9949 3224 16363 3226
rect 9949 3168 9954 3224
rect 10010 3168 16302 3224
rect 16358 3168 16363 3224
rect 9949 3166 16363 3168
rect 9949 3163 10015 3166
rect 16297 3163 16363 3166
rect 14733 3090 14799 3093
rect 16665 3090 16731 3093
rect 14733 3088 16731 3090
rect 14733 3032 14738 3088
rect 14794 3032 16670 3088
rect 16726 3032 16731 3088
rect 14733 3030 16731 3032
rect 14733 3027 14799 3030
rect 16665 3027 16731 3030
rect 16941 3090 17007 3093
rect 33501 3090 33567 3093
rect 16941 3088 33567 3090
rect 16941 3032 16946 3088
rect 17002 3032 33506 3088
rect 33562 3032 33567 3088
rect 16941 3030 33567 3032
rect 16941 3027 17007 3030
rect 33501 3027 33567 3030
rect 5165 2954 5231 2957
rect 19609 2954 19675 2957
rect 5165 2952 19675 2954
rect 5165 2896 5170 2952
rect 5226 2896 19614 2952
rect 19670 2896 19675 2952
rect 5165 2894 19675 2896
rect 5165 2891 5231 2894
rect 19609 2891 19675 2894
rect 15101 2818 15167 2821
rect 24577 2818 24643 2821
rect 15101 2816 24643 2818
rect 15101 2760 15106 2816
rect 15162 2760 24582 2816
rect 24638 2760 24643 2816
rect 15101 2758 24643 2760
rect 15101 2755 15167 2758
rect 24577 2755 24643 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 9949 2682 10015 2685
rect 13813 2682 13879 2685
rect 9949 2680 13879 2682
rect 9949 2624 9954 2680
rect 10010 2624 13818 2680
rect 13874 2624 13879 2680
rect 9949 2622 13879 2624
rect 9949 2619 10015 2622
rect 13813 2619 13879 2622
rect 16941 2546 17007 2549
rect 18638 2546 18644 2548
rect 16941 2544 18644 2546
rect 16941 2488 16946 2544
rect 17002 2488 18644 2544
rect 16941 2486 18644 2488
rect 16941 2483 17007 2486
rect 18638 2484 18644 2486
rect 18708 2484 18714 2548
rect 18781 2546 18847 2549
rect 37549 2546 37615 2549
rect 18781 2544 37615 2546
rect 18781 2488 18786 2544
rect 18842 2488 37554 2544
rect 37610 2488 37615 2544
rect 18781 2486 37615 2488
rect 18781 2483 18847 2486
rect 37549 2483 37615 2486
rect 4981 2410 5047 2413
rect 19609 2410 19675 2413
rect 4981 2408 19675 2410
rect 4981 2352 4986 2408
rect 5042 2352 19614 2408
rect 19670 2352 19675 2408
rect 4981 2350 19675 2352
rect 4981 2347 5047 2350
rect 19609 2347 19675 2350
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 9305 2002 9371 2005
rect 24209 2002 24275 2005
rect 9305 2000 24275 2002
rect 9305 1944 9310 2000
rect 9366 1944 24214 2000
rect 24270 1944 24275 2000
rect 9305 1942 24275 1944
rect 9305 1939 9371 1942
rect 24209 1939 24275 1942
rect 13077 1866 13143 1869
rect 27705 1866 27771 1869
rect 13077 1864 27771 1866
rect 13077 1808 13082 1864
rect 13138 1808 27710 1864
rect 27766 1808 27771 1864
rect 13077 1806 27771 1808
rect 13077 1803 13143 1806
rect 27705 1803 27771 1806
rect 19190 1668 19196 1732
rect 19260 1730 19266 1732
rect 31753 1730 31819 1733
rect 19260 1728 31819 1730
rect 19260 1672 31758 1728
rect 31814 1672 31819 1728
rect 19260 1670 31819 1672
rect 19260 1668 19266 1670
rect 31753 1667 31819 1670
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 21036 36484 21100 36548
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 36492 36000 36556 36004
rect 36492 35944 36542 36000
rect 36542 35944 36556 36000
rect 36492 35940 36556 35944
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 34652 34912 34716 34916
rect 34652 34856 34666 34912
rect 34666 34856 34716 34912
rect 34652 34852 34716 34856
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 23244 32948 23308 33012
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 36492 19952 36556 19956
rect 36492 19896 36506 19952
rect 36506 19896 36556 19952
rect 36492 19892 36556 19896
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 19380 17172 19444 17236
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 23244 15132 23308 15196
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 21036 14588 21100 14652
rect 34652 14588 34716 14652
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 18644 13832 18708 13836
rect 18644 13776 18694 13832
rect 18694 13776 18708 13832
rect 18644 13772 18708 13776
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19380 6836 19444 6900
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 19196 4116 19260 4180
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19380 3572 19444 3636
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 18644 2484 18708 2548
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 19196 1668 19260 1732
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 21035 36548 21101 36549
rect 21035 36484 21036 36548
rect 21100 36484 21101 36548
rect 21035 36483 21101 36484
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19379 17236 19445 17237
rect 19379 17172 19380 17236
rect 19444 17172 19445 17236
rect 19379 17171 19445 17172
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 18643 13836 18709 13837
rect 18643 13772 18644 13836
rect 18708 13772 18709 13836
rect 18643 13771 18709 13772
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 18646 2549 18706 13771
rect 19382 6901 19442 17171
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 21038 14653 21098 36483
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 36491 36004 36557 36005
rect 36491 35940 36492 36004
rect 36556 35940 36557 36004
rect 36491 35939 36557 35940
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34651 34916 34717 34917
rect 34651 34852 34652 34916
rect 34716 34852 34717 34916
rect 34651 34851 34717 34852
rect 23243 33012 23309 33013
rect 23243 32948 23244 33012
rect 23308 32948 23309 33012
rect 23243 32947 23309 32948
rect 23246 15197 23306 32947
rect 23243 15196 23309 15197
rect 23243 15132 23244 15196
rect 23308 15132 23309 15196
rect 23243 15131 23309 15132
rect 34654 14653 34714 34851
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 36494 19957 36554 35939
rect 36491 19956 36557 19957
rect 36491 19892 36492 19956
rect 36556 19892 36557 19956
rect 36491 19891 36557 19892
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 21035 14652 21101 14653
rect 21035 14588 21036 14652
rect 21100 14588 21101 14652
rect 21035 14587 21101 14588
rect 34651 14652 34717 14653
rect 34651 14588 34652 14652
rect 34716 14588 34717 14652
rect 34651 14587 34717 14588
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19379 6900 19445 6901
rect 19379 6836 19380 6900
rect 19444 6836 19445 6900
rect 19379 6835 19445 6836
rect 19195 4180 19261 4181
rect 19195 4116 19196 4180
rect 19260 4116 19261 4180
rect 19195 4115 19261 4116
rect 18643 2548 18709 2549
rect 18643 2484 18644 2548
rect 18708 2484 18709 2548
rect 18643 2483 18709 2484
rect 19198 1733 19258 4115
rect 19382 3637 19442 6835
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19379 3636 19445 3637
rect 19379 3572 19380 3636
rect 19444 3572 19445 3636
rect 19379 3571 19445 3572
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 19195 1732 19261 1733
rect 19195 1668 19196 1732
rect 19260 1668 19261 1732
rect 19195 1667 19261 1668
use sky130_fd_sc_hd__diode_2  ANTENNA__0438__A_N opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 37444 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0438__B
timestamp 1649977179
transform -1 0 37996 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0440__A
timestamp 1649977179
transform 1 0 15824 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0441__A
timestamp 1649977179
transform 1 0 16008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0442__B1
timestamp 1649977179
transform 1 0 16560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0443__A
timestamp 1649977179
transform 1 0 17664 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0447__A0
timestamp 1649977179
transform 1 0 18124 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0450__A0
timestamp 1649977179
transform 1 0 21804 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0452__A0
timestamp 1649977179
transform -1 0 19412 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0454__A0
timestamp 1649977179
transform 1 0 20884 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0456__A0
timestamp 1649977179
transform -1 0 21988 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__A0
timestamp 1649977179
transform 1 0 23000 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0460__A0
timestamp 1649977179
transform -1 0 21988 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0463__A0
timestamp 1649977179
transform 1 0 19596 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0465__A0
timestamp 1649977179
transform -1 0 23920 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0467__A0
timestamp 1649977179
transform 1 0 23184 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0469__A0
timestamp 1649977179
transform 1 0 25760 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0471__A0
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0473__A0
timestamp 1649977179
transform 1 0 22632 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0475__A0
timestamp 1649977179
transform 1 0 24196 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0477__A0
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0479__A0
timestamp 1649977179
transform 1 0 22632 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0481__A0
timestamp 1649977179
transform -1 0 19412 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0483__A0
timestamp 1649977179
transform 1 0 20976 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__A
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__B
timestamp 1649977179
transform 1 0 18216 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0489__A
timestamp 1649977179
transform -1 0 12420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0490__A
timestamp 1649977179
transform 1 0 18676 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0494__A
timestamp 1649977179
transform 1 0 17848 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__A
timestamp 1649977179
transform 1 0 19964 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__A2
timestamp 1649977179
transform 1 0 17112 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__A1
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__A2
timestamp 1649977179
transform -1 0 14628 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__A1
timestamp 1649977179
transform -1 0 14260 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__A2
timestamp 1649977179
transform -1 0 13616 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0503__A1
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0503__C1
timestamp 1649977179
transform 1 0 17480 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__A
timestamp 1649977179
transform 1 0 8740 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__B
timestamp 1649977179
transform 1 0 9752 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0507__A
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__A
timestamp 1649977179
transform 1 0 9476 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0510__A0
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0513__A
timestamp 1649977179
transform 1 0 15640 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0515__A
timestamp 1649977179
transform 1 0 13248 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0516__A1
timestamp 1649977179
transform 1 0 12328 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0518__B
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__C_N
timestamp 1649977179
transform 1 0 17020 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__A
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__B
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__A
timestamp 1649977179
transform 1 0 9108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__B
timestamp 1649977179
transform 1 0 9292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__A1
timestamp 1649977179
transform 1 0 14168 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__B1
timestamp 1649977179
transform 1 0 12512 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__A
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__A
timestamp 1649977179
transform 1 0 7728 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__B
timestamp 1649977179
transform 1 0 8280 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__A1
timestamp 1649977179
transform 1 0 8188 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__B
timestamp 1649977179
transform 1 0 16008 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__C_N
timestamp 1649977179
transform 1 0 15364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__A
timestamp 1649977179
transform -1 0 11776 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__B1
timestamp 1649977179
transform 1 0 15272 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0549__B
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__B1
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__A
timestamp 1649977179
transform 1 0 15824 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__B
timestamp 1649977179
transform 1 0 15272 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__A
timestamp 1649977179
transform -1 0 11132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__B
timestamp 1649977179
transform -1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0555__A
timestamp 1649977179
transform 1 0 28888 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0555__B
timestamp 1649977179
transform 1 0 29348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0557__A
timestamp 1649977179
transform 1 0 15364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__A
timestamp 1649977179
transform 1 0 31832 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__B
timestamp 1649977179
transform 1 0 31464 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__A1
timestamp 1649977179
transform 1 0 23184 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__B1
timestamp 1649977179
transform 1 0 22356 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0563__A1
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__A1
timestamp 1649977179
transform -1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__A2
timestamp 1649977179
transform 1 0 19872 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__A0
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__A1
timestamp 1649977179
transform -1 0 20240 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__S
timestamp 1649977179
transform 1 0 18584 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__A0
timestamp 1649977179
transform -1 0 21160 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__A1
timestamp 1649977179
transform 1 0 20424 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__S
timestamp 1649977179
transform 1 0 18584 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__S
timestamp 1649977179
transform 1 0 35604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__S
timestamp 1649977179
transform 1 0 35972 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__A0
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__S
timestamp 1649977179
transform -1 0 33120 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__A1
timestamp 1649977179
transform -1 0 12328 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__S
timestamp 1649977179
transform -1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__A1
timestamp 1649977179
transform -1 0 15272 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__S
timestamp 1649977179
transform 1 0 14812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__A1
timestamp 1649977179
transform -1 0 16836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__S
timestamp 1649977179
transform 1 0 15824 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__A1
timestamp 1649977179
transform -1 0 33212 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__S
timestamp 1649977179
transform 1 0 33580 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__A1
timestamp 1649977179
transform -1 0 31556 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__S
timestamp 1649977179
transform 1 0 31464 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__S
timestamp 1649977179
transform 1 0 29900 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__A1
timestamp 1649977179
transform -1 0 33488 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__S
timestamp 1649977179
transform 1 0 31924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A1
timestamp 1649977179
transform -1 0 37996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__S
timestamp 1649977179
transform 1 0 33212 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__A1
timestamp 1649977179
transform 1 0 31464 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__S
timestamp 1649977179
transform 1 0 30544 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__A1
timestamp 1649977179
transform 1 0 36616 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__S
timestamp 1649977179
transform 1 0 32476 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__A1
timestamp 1649977179
transform 1 0 35696 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__S
timestamp 1649977179
transform -1 0 33396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__A1
timestamp 1649977179
transform 1 0 36248 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__S
timestamp 1649977179
transform -1 0 35328 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__A1
timestamp 1649977179
transform 1 0 36340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__S
timestamp 1649977179
transform -1 0 36524 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__S
timestamp 1649977179
transform -1 0 34776 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__A1
timestamp 1649977179
transform -1 0 35972 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__S
timestamp 1649977179
transform 1 0 35236 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__A1
timestamp 1649977179
transform -1 0 35420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__S
timestamp 1649977179
transform 1 0 33488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__A1
timestamp 1649977179
transform -1 0 23644 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__S
timestamp 1649977179
transform -1 0 17756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__A1
timestamp 1649977179
transform -1 0 20608 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__S
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A1
timestamp 1649977179
transform -1 0 23092 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__S
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A1
timestamp 1649977179
transform -1 0 12880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A1
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__A1
timestamp 1649977179
transform 1 0 11040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__A1
timestamp 1649977179
transform 1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__A1
timestamp 1649977179
transform -1 0 6256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__A1
timestamp 1649977179
transform -1 0 12696 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__A1
timestamp 1649977179
transform -1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__A1
timestamp 1649977179
transform -1 0 8740 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A1
timestamp 1649977179
transform -1 0 7268 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__A1
timestamp 1649977179
transform -1 0 8464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__A1
timestamp 1649977179
transform -1 0 16836 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A1
timestamp 1649977179
transform 1 0 15364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__A1
timestamp 1649977179
transform -1 0 15272 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__A1
timestamp 1649977179
transform 1 0 14720 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__A1
timestamp 1649977179
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__A1
timestamp 1649977179
transform -1 0 18032 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A1
timestamp 1649977179
transform 1 0 18584 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__A1
timestamp 1649977179
transform -1 0 20332 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__A1
timestamp 1649977179
transform -1 0 18584 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__A1
timestamp 1649977179
transform 1 0 20884 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__A1
timestamp 1649977179
transform -1 0 20240 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__A1
timestamp 1649977179
transform 1 0 17296 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__A
timestamp 1649977179
transform 1 0 15732 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A0
timestamp 1649977179
transform 1 0 18032 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A1
timestamp 1649977179
transform -1 0 18584 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A
timestamp 1649977179
transform 1 0 15456 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A0
timestamp 1649977179
transform 1 0 18584 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A1
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__A
timestamp 1649977179
transform 1 0 16008 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A0
timestamp 1649977179
transform -1 0 17296 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A1
timestamp 1649977179
transform 1 0 18216 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A
timestamp 1649977179
transform -1 0 14996 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A0
timestamp 1649977179
transform -1 0 19688 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A1
timestamp 1649977179
transform 1 0 18952 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A
timestamp 1649977179
transform 1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A0
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A1
timestamp 1649977179
transform 1 0 22264 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A1
timestamp 1649977179
transform -1 0 22816 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A
timestamp 1649977179
transform 1 0 17664 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A0
timestamp 1649977179
transform -1 0 19780 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A1
timestamp 1649977179
transform -1 0 20148 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A
timestamp 1649977179
transform 1 0 20056 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A0
timestamp 1649977179
transform 1 0 20976 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A1
timestamp 1649977179
transform -1 0 20608 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A
timestamp 1649977179
transform 1 0 18216 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A0
timestamp 1649977179
transform -1 0 22356 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A1
timestamp 1649977179
transform -1 0 21252 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A0
timestamp 1649977179
transform 1 0 20792 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A1
timestamp 1649977179
transform 1 0 21160 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__A0
timestamp 1649977179
transform -1 0 23092 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__A1
timestamp 1649977179
transform 1 0 23460 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A0
timestamp 1649977179
transform -1 0 21068 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A1
timestamp 1649977179
transform -1 0 21988 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A0
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A1
timestamp 1649977179
transform 1 0 22724 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A0
timestamp 1649977179
transform 1 0 23920 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A1
timestamp 1649977179
transform -1 0 24656 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A0
timestamp 1649977179
transform -1 0 25484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A1
timestamp 1649977179
transform -1 0 25944 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A0
timestamp 1649977179
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A1
timestamp 1649977179
transform 1 0 26312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A0
timestamp 1649977179
transform 1 0 26312 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A1
timestamp 1649977179
transform -1 0 27140 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A
timestamp 1649977179
transform -1 0 24472 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B
timestamp 1649977179
transform -1 0 24012 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__A
timestamp 1649977179
transform -1 0 32292 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 1649977179
transform 1 0 30176 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1649977179
transform -1 0 17848 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__B
timestamp 1649977179
transform 1 0 16008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A
timestamp 1649977179
transform -1 0 17112 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A0
timestamp 1649977179
transform -1 0 26772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A1
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__S
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A
timestamp 1649977179
transform -1 0 24564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A0
timestamp 1649977179
transform 1 0 24932 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A1
timestamp 1649977179
transform -1 0 23920 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__S
timestamp 1649977179
transform 1 0 23276 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A
timestamp 1649977179
transform 1 0 23092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A0
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A1
timestamp 1649977179
transform -1 0 21896 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__S
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A
timestamp 1649977179
transform 1 0 22724 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A0
timestamp 1649977179
transform -1 0 36524 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__S
timestamp 1649977179
transform 1 0 34960 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A
timestamp 1649977179
transform 1 0 28888 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__S
timestamp 1649977179
transform 1 0 35512 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__S
timestamp 1649977179
transform -1 0 36800 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A0
timestamp 1649977179
transform -1 0 23368 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A1
timestamp 1649977179
transform 1 0 22632 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__S
timestamp 1649977179
transform 1 0 21620 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A0
timestamp 1649977179
transform -1 0 27324 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A1
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__S
timestamp 1649977179
transform 1 0 25576 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A0
timestamp 1649977179
transform -1 0 30268 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A1
timestamp 1649977179
transform -1 0 29716 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__S
timestamp 1649977179
transform 1 0 27784 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A0
timestamp 1649977179
transform -1 0 30360 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A1
timestamp 1649977179
transform 1 0 29624 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__S
timestamp 1649977179
transform 1 0 29072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A0
timestamp 1649977179
transform -1 0 28428 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A1
timestamp 1649977179
transform 1 0 28796 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A0
timestamp 1649977179
transform -1 0 30544 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A1
timestamp 1649977179
transform -1 0 32292 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A0
timestamp 1649977179
transform -1 0 31464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A1
timestamp 1649977179
transform 1 0 30728 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A
timestamp 1649977179
transform 1 0 18768 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A0
timestamp 1649977179
transform -1 0 32844 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A1
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A
timestamp 1649977179
transform -1 0 30820 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A0
timestamp 1649977179
transform 1 0 34684 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A1
timestamp 1649977179
transform 1 0 34224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A
timestamp 1649977179
transform 1 0 32384 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A0
timestamp 1649977179
transform -1 0 37076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A1
timestamp 1649977179
transform -1 0 35328 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A
timestamp 1649977179
transform -1 0 36340 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A1
timestamp 1649977179
transform 1 0 35512 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A
timestamp 1649977179
transform -1 0 33488 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A1
timestamp 1649977179
transform -1 0 37260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A
timestamp 1649977179
transform 1 0 35788 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A
timestamp 1649977179
transform 1 0 35236 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A0
timestamp 1649977179
transform 1 0 34224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A1
timestamp 1649977179
transform -1 0 33856 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__S
timestamp 1649977179
transform 1 0 33948 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A
timestamp 1649977179
transform 1 0 33304 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A1
timestamp 1649977179
transform 1 0 36340 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__S
timestamp 1649977179
transform 1 0 33856 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A
timestamp 1649977179
transform -1 0 37168 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A0
timestamp 1649977179
transform 1 0 20424 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A1
timestamp 1649977179
transform 1 0 19780 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__S
timestamp 1649977179
transform 1 0 19964 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A
timestamp 1649977179
transform -1 0 19596 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A0
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A1
timestamp 1649977179
transform -1 0 18492 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__S
timestamp 1649977179
transform 1 0 16836 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A
timestamp 1649977179
transform 1 0 18400 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A
timestamp 1649977179
transform -1 0 13800 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A0
timestamp 1649977179
transform 1 0 15272 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A1
timestamp 1649977179
transform 1 0 15824 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__S
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A0
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A1
timestamp 1649977179
transform -1 0 11684 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__S
timestamp 1649977179
transform 1 0 12788 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A0
timestamp 1649977179
transform 1 0 10212 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A1
timestamp 1649977179
transform -1 0 10948 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__S
timestamp 1649977179
transform -1 0 9844 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A0
timestamp 1649977179
transform 1 0 10120 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A1
timestamp 1649977179
transform -1 0 10856 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__S
timestamp 1649977179
transform 1 0 9752 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A0
timestamp 1649977179
transform 1 0 10304 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A1
timestamp 1649977179
transform 1 0 10120 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__S
timestamp 1649977179
transform 1 0 10672 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A0
timestamp 1649977179
transform -1 0 12880 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A1
timestamp 1649977179
transform 1 0 12512 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__S
timestamp 1649977179
transform 1 0 12788 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A0
timestamp 1649977179
transform -1 0 13708 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A1
timestamp 1649977179
transform 1 0 13156 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__A0
timestamp 1649977179
transform 1 0 13432 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__A1
timestamp 1649977179
transform -1 0 13248 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A0
timestamp 1649977179
transform 1 0 13156 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A1
timestamp 1649977179
transform -1 0 13708 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A0
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A1
timestamp 1649977179
transform -1 0 12604 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A
timestamp 1649977179
transform 1 0 15640 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A0
timestamp 1649977179
transform -1 0 14444 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A1
timestamp 1649977179
transform -1 0 14260 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A0
timestamp 1649977179
transform 1 0 16376 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A1
timestamp 1649977179
transform 1 0 16008 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A0
timestamp 1649977179
transform -1 0 16560 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A1
timestamp 1649977179
transform -1 0 16376 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__A0
timestamp 1649977179
transform -1 0 15824 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__A1
timestamp 1649977179
transform 1 0 15272 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A0
timestamp 1649977179
transform -1 0 16836 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A1
timestamp 1649977179
transform -1 0 15640 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A0
timestamp 1649977179
transform -1 0 16192 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A1
timestamp 1649977179
transform -1 0 16376 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A0
timestamp 1649977179
transform -1 0 17940 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A1
timestamp 1649977179
transform 1 0 17204 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A0
timestamp 1649977179
transform -1 0 18032 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A1
timestamp 1649977179
transform 1 0 17480 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A0
timestamp 1649977179
transform 1 0 18216 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A1
timestamp 1649977179
transform -1 0 16652 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A0
timestamp 1649977179
transform 1 0 20424 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A0
timestamp 1649977179
transform 1 0 22908 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A1
timestamp 1649977179
transform -1 0 22540 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A
timestamp 1649977179
transform 1 0 19780 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A0
timestamp 1649977179
transform 1 0 21068 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A1
timestamp 1649977179
transform -1 0 20700 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A
timestamp 1649977179
transform 1 0 20148 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A0
timestamp 1649977179
transform 1 0 22172 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A1
timestamp 1649977179
transform -1 0 21344 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A
timestamp 1649977179
transform 1 0 22632 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__D
timestamp 1649977179
transform -1 0 29072 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__D
timestamp 1649977179
transform -1 0 30820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__D
timestamp 1649977179
transform 1 0 28888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__D
timestamp 1649977179
transform -1 0 37444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__D
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__D
timestamp 1649977179
transform -1 0 35420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__D
timestamp 1649977179
transform -1 0 30912 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_m_A
timestamp 1649977179
transform -1 0 32292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_s_A
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 1840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 2392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 4048 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 5704 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 7912 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 6716 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 6808 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 7820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 8924 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 5244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 9476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 7360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 4784 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 14444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 11684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 10028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 5428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 6072 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 5336 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 5152 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 5888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 7636 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 8004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 6808 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 11224 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 29716 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 34040 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 38180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 35972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 37444 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 37904 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 37444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 29532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 29072 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 30084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 31556 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 30636 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 33948 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 32936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 31648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 37628 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 38180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 37996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 37996 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 38180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 2024 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 3128 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 17020 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 17940 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 26220 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 23920 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 25116 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 27784 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 28060 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 27508 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 17572 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 18584 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 18124 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 26496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 20976 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 23368 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 26312 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 29716 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output68_A
timestamp 1649977179
transform -1 0 3128 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output69_A
timestamp 1649977179
transform -1 0 11684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output70_A
timestamp 1649977179
transform 1 0 25944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output71_A
timestamp 1649977179
transform 1 0 28888 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1649977179
transform 1 0 25576 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output73_A
timestamp 1649977179
transform 1 0 31464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output74_A
timestamp 1649977179
transform 1 0 30084 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output75_A
timestamp 1649977179
transform 1 0 28796 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1649977179
transform 1 0 19412 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output77_A
timestamp 1649977179
transform -1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output78_A
timestamp 1649977179
transform 1 0 21160 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output80_A
timestamp 1649977179
transform 1 0 22356 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output81_A
timestamp 1649977179
transform 1 0 24748 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output82_A
timestamp 1649977179
transform -1 0 26496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output83_A
timestamp 1649977179
transform 1 0 23552 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output84_A
timestamp 1649977179
transform 1 0 26128 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output85_A
timestamp 1649977179
transform 1 0 2576 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1649977179
transform -1 0 2576 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output87_A
timestamp 1649977179
transform 1 0 4416 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1649977179
transform 1 0 9568 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output89_A
timestamp 1649977179
transform 1 0 10304 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output90_A
timestamp 1649977179
transform 1 0 11040 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output91_A
timestamp 1649977179
transform -1 0 10304 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output92_A
timestamp 1649977179
transform 1 0 12144 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output93_A
timestamp 1649977179
transform 1 0 12696 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1649977179
transform -1 0 11960 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output95_A
timestamp 1649977179
transform 1 0 13432 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output96_A
timestamp 1649977179
transform 1 0 14352 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output97_A
timestamp 1649977179
transform -1 0 13616 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output98_A
timestamp 1649977179
transform 1 0 4968 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output99_A
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output100_A
timestamp 1649977179
transform -1 0 15272 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output101_A
timestamp 1649977179
transform -1 0 15916 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output102_A
timestamp 1649977179
transform 1 0 17112 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output103_A
timestamp 1649977179
transform 1 0 5520 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output104_A
timestamp 1649977179
transform 1 0 5704 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output105_A
timestamp 1649977179
transform 1 0 6716 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output106_A
timestamp 1649977179
transform 1 0 7268 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output107_A
timestamp 1649977179
transform 1 0 7360 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output108_A
timestamp 1649977179
transform 1 0 8280 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output109_A
timestamp 1649977179
transform 1 0 8464 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output110_A
timestamp 1649977179
transform 1 0 9384 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output111_A
timestamp 1649977179
transform -1 0 16468 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output112_A
timestamp 1649977179
transform 1 0 28428 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output113_A
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output117_A
timestamp 1649977179
transform -1 0 38180 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 1649977179
transform 1 0 29992 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output120_A
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output121_A
timestamp 1649977179
transform 1 0 30544 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output122_A
timestamp 1649977179
transform 1 0 31096 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output123_A
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output125_A
timestamp 1649977179
transform -1 0 34868 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output126_A
timestamp 1649977179
transform 1 0 34960 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output127_A
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output128_A
timestamp 1649977179
transform -1 0 35696 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39
timestamp 1649977179
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1649977179
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1649977179
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1649977179
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1649977179
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115
timestamp 1649977179
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122
timestamp 1649977179
transform 1 0 12328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_143
timestamp 1649977179
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150
timestamp 1649977179
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_176
timestamp 1649977179
transform 1 0 17296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1649977179
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1649977179
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1649977179
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1649977179
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_229
timestamp 1649977179
transform 1 0 22172 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1649977179
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1649977179
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1649977179
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_285
timestamp 1649977179
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_293
timestamp 1649977179
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1649977179
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_312
timestamp 1649977179
transform 1 0 29808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_319
timestamp 1649977179
transform 1 0 30452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_326
timestamp 1649977179
transform 1 0 31096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1649977179
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_341
timestamp 1649977179
transform 1 0 32476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_358
timestamp 1649977179
transform 1 0 34040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1649977179
transform 1 0 34960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1649977179
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_8
timestamp 1649977179
transform 1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_14
timestamp 1649977179
transform 1 0 2392 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1649977179
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1649977179
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_34
timestamp 1649977179
transform 1 0 4232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1649977179
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1649977179
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_61
timestamp 1649977179
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_65
timestamp 1649977179
transform 1 0 7084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1649977179
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_80
timestamp 1649977179
transform 1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_104 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10672 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_123
timestamp 1649977179
transform 1 0 12420 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1649977179
transform 1 0 13248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1649977179
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_145
timestamp 1649977179
transform 1 0 14444 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1649977179
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_189
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_206
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp 1649977179
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_241
timestamp 1649977179
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_249
timestamp 1649977179
transform 1 0 24012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_253
timestamp 1649977179
transform 1 0 24380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_270
timestamp 1649977179
transform 1 0 25944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1649977179
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_324
timestamp 1649977179
transform 1 0 30912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_328
timestamp 1649977179
transform 1 0 31280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1649977179
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_353
timestamp 1649977179
transform 1 0 33580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_360
timestamp 1649977179
transform 1 0 34224 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_368
timestamp 1649977179
transform 1 0 34960 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1649977179
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_393
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1649977179
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_21
timestamp 1649977179
transform 1 0 3036 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_35
timestamp 1649977179
transform 1 0 4324 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_44
timestamp 1649977179
transform 1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_50
timestamp 1649977179
transform 1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_56
timestamp 1649977179
transform 1 0 6256 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_62
timestamp 1649977179
transform 1 0 6808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1649977179
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_74
timestamp 1649977179
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_90
timestamp 1649977179
transform 1 0 9384 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_101
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_105
timestamp 1649977179
transform 1 0 10764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_116
timestamp 1649977179
transform 1 0 11776 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1649977179
transform 1 0 12880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_132
timestamp 1649977179
transform 1 0 13248 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1649977179
transform 1 0 14720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_156
timestamp 1649977179
transform 1 0 15456 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_170
timestamp 1649977179
transform 1 0 16744 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_178
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_206
timestamp 1649977179
transform 1 0 20056 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_214
timestamp 1649977179
transform 1 0 20792 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_236
timestamp 1649977179
transform 1 0 22816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_244
timestamp 1649977179
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_257
timestamp 1649977179
transform 1 0 24748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_291
timestamp 1649977179
transform 1 0 27876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_298
timestamp 1649977179
transform 1 0 28520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1649977179
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_311
timestamp 1649977179
transform 1 0 29716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_317
timestamp 1649977179
transform 1 0 30268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_323
timestamp 1649977179
transform 1 0 30820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_347
timestamp 1649977179
transform 1 0 33028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1649977179
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_384
timestamp 1649977179
transform 1 0 36432 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_391
timestamp 1649977179
transform 1 0 37076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_398
timestamp 1649977179
transform 1 0 37720 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_406
timestamp 1649977179
transform 1 0 38456 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_32
timestamp 1649977179
transform 1 0 4048 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_40
timestamp 1649977179
transform 1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_46
timestamp 1649977179
transform 1 0 5336 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_61
timestamp 1649977179
transform 1 0 6716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_67
timestamp 1649977179
transform 1 0 7268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_73
timestamp 1649977179
transform 1 0 7820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_79
timestamp 1649977179
transform 1 0 8372 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1649977179
transform 1 0 8924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_91
timestamp 1649977179
transform 1 0 9476 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1649977179
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1649977179
transform 1 0 11684 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_122
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_129
timestamp 1649977179
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_136
timestamp 1649977179
transform 1 0 13616 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_143
timestamp 1649977179
transform 1 0 14260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_151
timestamp 1649977179
transform 1 0 14996 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_154
timestamp 1649977179
transform 1 0 15272 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_171
timestamp 1649977179
transform 1 0 16836 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_192
timestamp 1649977179
transform 1 0 18768 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1649977179
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_214
timestamp 1649977179
transform 1 0 20792 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_227
timestamp 1649977179
transform 1 0 21988 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_233
timestamp 1649977179
transform 1 0 22540 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_239
timestamp 1649977179
transform 1 0 23092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_245
timestamp 1649977179
transform 1 0 23644 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_266
timestamp 1649977179
transform 1 0 25576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_272
timestamp 1649977179
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_298
timestamp 1649977179
transform 1 0 28520 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_325
timestamp 1649977179
transform 1 0 31004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp 1649977179
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_346
timestamp 1649977179
transform 1 0 32936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_350
timestamp 1649977179
transform 1 0 33304 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_360
timestamp 1649977179
transform 1 0 34224 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_367
timestamp 1649977179
transform 1 0 34868 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_371
timestamp 1649977179
transform 1 0 35236 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1649977179
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_396
timestamp 1649977179
transform 1 0 37536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1649977179
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_47
timestamp 1649977179
transform 1 0 5428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_51
timestamp 1649977179
transform 1 0 5796 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_54
timestamp 1649977179
transform 1 0 6072 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_62
timestamp 1649977179
transform 1 0 6808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_68
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_74
timestamp 1649977179
transform 1 0 7912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_91
timestamp 1649977179
transform 1 0 9476 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_104
timestamp 1649977179
transform 1 0 10672 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_110
timestamp 1649977179
transform 1 0 11224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_116
timestamp 1649977179
transform 1 0 11776 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_122
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_131
timestamp 1649977179
transform 1 0 13156 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_146
timestamp 1649977179
transform 1 0 14536 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_156
timestamp 1649977179
transform 1 0 15456 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_162
timestamp 1649977179
transform 1 0 16008 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_169
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_175
timestamp 1649977179
transform 1 0 17204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_181
timestamp 1649977179
transform 1 0 17756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_188
timestamp 1649977179
transform 1 0 18400 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_203
timestamp 1649977179
transform 1 0 19780 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_211
timestamp 1649977179
transform 1 0 20516 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_217
timestamp 1649977179
transform 1 0 21068 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_239
timestamp 1649977179
transform 1 0 23092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_243
timestamp 1649977179
transform 1 0 23460 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_246
timestamp 1649977179
transform 1 0 23736 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_258
timestamp 1649977179
transform 1 0 24840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_278
timestamp 1649977179
transform 1 0 26680 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_298
timestamp 1649977179
transform 1 0 28520 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1649977179
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_316
timestamp 1649977179
transform 1 0 30176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_322
timestamp 1649977179
transform 1 0 30728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_335
timestamp 1649977179
transform 1 0 31924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_342
timestamp 1649977179
transform 1 0 32568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_349
timestamp 1649977179
transform 1 0 33212 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1649977179
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_374
timestamp 1649977179
transform 1 0 35512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_378
timestamp 1649977179
transform 1 0 35880 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_395
timestamp 1649977179
transform 1 0 37444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_399
timestamp 1649977179
transform 1 0 37812 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1649977179
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_71
timestamp 1649977179
transform 1 0 7636 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_77
timestamp 1649977179
transform 1 0 8188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_83
timestamp 1649977179
transform 1 0 8740 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_89
timestamp 1649977179
transform 1 0 9292 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_95
timestamp 1649977179
transform 1 0 9844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_118
timestamp 1649977179
transform 1 0 11960 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_124
timestamp 1649977179
transform 1 0 12512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_131
timestamp 1649977179
transform 1 0 13156 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_143
timestamp 1649977179
transform 1 0 14260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_153
timestamp 1649977179
transform 1 0 15180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_175
timestamp 1649977179
transform 1 0 17204 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_183
timestamp 1649977179
transform 1 0 17940 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_187
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_196
timestamp 1649977179
transform 1 0 19136 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_204
timestamp 1649977179
transform 1 0 19872 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_210
timestamp 1649977179
transform 1 0 20424 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_227
timestamp 1649977179
transform 1 0 21988 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_239
timestamp 1649977179
transform 1 0 23092 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_262
timestamp 1649977179
transform 1 0 25208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_268
timestamp 1649977179
transform 1 0 25760 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1649977179
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_297
timestamp 1649977179
transform 1 0 28428 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_303
timestamp 1649977179
transform 1 0 28980 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_309
timestamp 1649977179
transform 1 0 29532 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_315
timestamp 1649977179
transform 1 0 30084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_321
timestamp 1649977179
transform 1 0 30636 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1649977179
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_350
timestamp 1649977179
transform 1 0 33304 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_354
timestamp 1649977179
transform 1 0 33672 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_375
timestamp 1649977179
transform 1 0 35604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_382
timestamp 1649977179
transform 1 0 36248 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1649977179
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_396
timestamp 1649977179
transform 1 0 37536 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1649977179
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1649977179
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_105
timestamp 1649977179
transform 1 0 10764 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_115
timestamp 1649977179
transform 1 0 11684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_129
timestamp 1649977179
transform 1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_145
timestamp 1649977179
transform 1 0 14444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_151
timestamp 1649977179
transform 1 0 14996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_157
timestamp 1649977179
transform 1 0 15548 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_161
timestamp 1649977179
transform 1 0 15916 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_164
timestamp 1649977179
transform 1 0 16192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_186
timestamp 1649977179
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1649977179
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_207
timestamp 1649977179
transform 1 0 20148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1649977179
transform 1 0 20884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_222
timestamp 1649977179
transform 1 0 21528 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_244
timestamp 1649977179
transform 1 0 23552 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_259
timestamp 1649977179
transform 1 0 24932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_271
timestamp 1649977179
transform 1 0 26036 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_279
timestamp 1649977179
transform 1 0 26772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_296
timestamp 1649977179
transform 1 0 28336 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1649977179
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_325
timestamp 1649977179
transform 1 0 31004 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_331
timestamp 1649977179
transform 1 0 31556 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_337
timestamp 1649977179
transform 1 0 32108 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_343
timestamp 1649977179
transform 1 0 32660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_349
timestamp 1649977179
transform 1 0 33212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_355
timestamp 1649977179
transform 1 0 33764 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_374
timestamp 1649977179
transform 1 0 35512 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_378
timestamp 1649977179
transform 1 0 35880 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_382
timestamp 1649977179
transform 1 0 36248 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_386
timestamp 1649977179
transform 1 0 36616 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1649977179
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1649977179
transform 1 0 10120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_122
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_129
timestamp 1649977179
transform 1 0 12972 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_140
timestamp 1649977179
transform 1 0 13984 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_146
timestamp 1649977179
transform 1 0 14536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1649977179
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1649977179
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_176
timestamp 1649977179
transform 1 0 17296 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_182
timestamp 1649977179
transform 1 0 17848 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_189
timestamp 1649977179
transform 1 0 18492 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_195
timestamp 1649977179
transform 1 0 19044 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_201
timestamp 1649977179
transform 1 0 19596 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_208
timestamp 1649977179
transform 1 0 20240 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_216
timestamp 1649977179
transform 1 0 20976 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1649977179
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_241
timestamp 1649977179
transform 1 0 23276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_253
timestamp 1649977179
transform 1 0 24380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_270
timestamp 1649977179
transform 1 0 25944 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1649977179
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_313
timestamp 1649977179
transform 1 0 29900 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_326
timestamp 1649977179
transform 1 0 31096 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1649977179
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_346
timestamp 1649977179
transform 1 0 32936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_352
timestamp 1649977179
transform 1 0 33488 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_358
timestamp 1649977179
transform 1 0 34040 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_367
timestamp 1649977179
transform 1 0 34868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_379
timestamp 1649977179
transform 1 0 35972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_398
timestamp 1649977179
transform 1 0 37720 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_406
timestamp 1649977179
transform 1 0 38456 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_105
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_116
timestamp 1649977179
transform 1 0 11776 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_126
timestamp 1649977179
transform 1 0 12696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_148
timestamp 1649977179
transform 1 0 14720 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_156
timestamp 1649977179
transform 1 0 15456 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_162
timestamp 1649977179
transform 1 0 16008 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_171
timestamp 1649977179
transform 1 0 16836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_178
timestamp 1649977179
transform 1 0 17480 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_184
timestamp 1649977179
transform 1 0 18032 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_206
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_213
timestamp 1649977179
transform 1 0 20700 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_239
timestamp 1649977179
transform 1 0 23092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_284
timestamp 1649977179
transform 1 0 27232 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_296
timestamp 1649977179
transform 1 0 28336 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_315
timestamp 1649977179
transform 1 0 30084 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_328
timestamp 1649977179
transform 1 0 31280 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_348
timestamp 1649977179
transform 1 0 33120 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_356
timestamp 1649977179
transform 1 0 33856 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1649977179
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_374
timestamp 1649977179
transform 1 0 35512 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_380
timestamp 1649977179
transform 1 0 36064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_397
timestamp 1649977179
transform 1 0 37628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_403
timestamp 1649977179
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_89
timestamp 1649977179
transform 1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_95
timestamp 1649977179
transform 1 0 9844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_120
timestamp 1649977179
transform 1 0 12144 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_128
timestamp 1649977179
transform 1 0 12880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_131
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_138
timestamp 1649977179
transform 1 0 13800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_144
timestamp 1649977179
transform 1 0 14352 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_152
timestamp 1649977179
transform 1 0 15088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_158
timestamp 1649977179
transform 1 0 15640 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1649977179
transform 1 0 17848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_192
timestamp 1649977179
transform 1 0 18768 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_198
timestamp 1649977179
transform 1 0 19320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_202
timestamp 1649977179
transform 1 0 19688 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_208
timestamp 1649977179
transform 1 0 20240 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1649977179
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1649977179
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_301
timestamp 1649977179
transform 1 0 28796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_325
timestamp 1649977179
transform 1 0 31004 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp 1649977179
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_340
timestamp 1649977179
transform 1 0 32384 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_346
timestamp 1649977179
transform 1 0 32936 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_354
timestamp 1649977179
transform 1 0 33672 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_367
timestamp 1649977179
transform 1 0 34868 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_379
timestamp 1649977179
transform 1 0 35972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_395
timestamp 1649977179
transform 1 0 37444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_401
timestamp 1649977179
transform 1 0 37996 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_105
timestamp 1649977179
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_110
timestamp 1649977179
transform 1 0 11224 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_122
timestamp 1649977179
transform 1 0 12328 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_126
timestamp 1649977179
transform 1 0 12696 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_149
timestamp 1649977179
transform 1 0 14812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_164
timestamp 1649977179
transform 1 0 16192 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_170
timestamp 1649977179
transform 1 0 16744 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_185
timestamp 1649977179
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1649977179
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_200
timestamp 1649977179
transform 1 0 19504 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_206
timestamp 1649977179
transform 1 0 20056 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_218
timestamp 1649977179
transform 1 0 21160 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_240
timestamp 1649977179
transform 1 0 23184 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_315
timestamp 1649977179
transform 1 0 30084 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_336
timestamp 1649977179
transform 1 0 32016 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_356
timestamp 1649977179
transform 1 0 33856 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_374
timestamp 1649977179
transform 1 0 35512 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_383
timestamp 1649977179
transform 1 0 36340 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_403
timestamp 1649977179
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_101
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1649977179
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_124
timestamp 1649977179
transform 1 0 12512 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_130
timestamp 1649977179
transform 1 0 13064 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_138
timestamp 1649977179
transform 1 0 13800 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_148
timestamp 1649977179
transform 1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_152
timestamp 1649977179
transform 1 0 15088 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_156
timestamp 1649977179
transform 1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_162
timestamp 1649977179
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_175
timestamp 1649977179
transform 1 0 17204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_198
timestamp 1649977179
transform 1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_202
timestamp 1649977179
transform 1 0 19688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_211
timestamp 1649977179
transform 1 0 20516 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_241
timestamp 1649977179
transform 1 0 23276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_253
timestamp 1649977179
transform 1 0 24380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_265
timestamp 1649977179
transform 1 0 25484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1649977179
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_297
timestamp 1649977179
transform 1 0 28428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_309
timestamp 1649977179
transform 1 0 29532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_321
timestamp 1649977179
transform 1 0 30636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 1649977179
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_339
timestamp 1649977179
transform 1 0 32292 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_347
timestamp 1649977179
transform 1 0 33028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_351
timestamp 1649977179
transform 1 0 33396 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_360
timestamp 1649977179
transform 1 0 34224 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_366
timestamp 1649977179
transform 1 0 34776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_372
timestamp 1649977179
transform 1 0 35328 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_378
timestamp 1649977179
transform 1 0 35880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_384
timestamp 1649977179
transform 1 0 36432 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_395
timestamp 1649977179
transform 1 0 37444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_401
timestamp 1649977179
transform 1 0 37996 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_93
timestamp 1649977179
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_105
timestamp 1649977179
transform 1 0 10764 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_113
timestamp 1649977179
transform 1 0 11500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_117
timestamp 1649977179
transform 1 0 11868 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_123
timestamp 1649977179
transform 1 0 12420 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_144
timestamp 1649977179
transform 1 0 14352 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_150
timestamp 1649977179
transform 1 0 14904 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_162
timestamp 1649977179
transform 1 0 16008 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_170
timestamp 1649977179
transform 1 0 16744 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_174
timestamp 1649977179
transform 1 0 17112 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_181
timestamp 1649977179
transform 1 0 17756 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1649977179
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_206
timestamp 1649977179
transform 1 0 20056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_212
timestamp 1649977179
transform 1 0 20608 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1649977179
transform 1 0 21160 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_238
timestamp 1649977179
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1649977179
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_259
timestamp 1649977179
transform 1 0 24932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_276
timestamp 1649977179
transform 1 0 26496 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_284
timestamp 1649977179
transform 1 0 27232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_302
timestamp 1649977179
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_317
timestamp 1649977179
transform 1 0 30268 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_336
timestamp 1649977179
transform 1 0 32016 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_348
timestamp 1649977179
transform 1 0 33120 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_351
timestamp 1649977179
transform 1 0 33396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_368
timestamp 1649977179
transform 1 0 34960 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_374
timestamp 1649977179
transform 1 0 35512 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_391
timestamp 1649977179
transform 1 0 37076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_397
timestamp 1649977179
transform 1 0 37628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1649977179
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1649977179
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_122
timestamp 1649977179
transform 1 0 12328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_128
timestamp 1649977179
transform 1 0 12880 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_136
timestamp 1649977179
transform 1 0 13616 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_148
timestamp 1649977179
transform 1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_154
timestamp 1649977179
transform 1 0 15272 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1649977179
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_176
timestamp 1649977179
transform 1 0 17296 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_182
timestamp 1649977179
transform 1 0 17848 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_190
timestamp 1649977179
transform 1 0 18584 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_194
timestamp 1649977179
transform 1 0 18952 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_200
timestamp 1649977179
transform 1 0 19504 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_209
timestamp 1649977179
transform 1 0 20332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_216
timestamp 1649977179
transform 1 0 20976 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_245
timestamp 1649977179
transform 1 0 23644 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_265
timestamp 1649977179
transform 1 0 25484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1649977179
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_297
timestamp 1649977179
transform 1 0 28428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_322
timestamp 1649977179
transform 1 0 30728 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1649977179
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_345
timestamp 1649977179
transform 1 0 32844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_363
timestamp 1649977179
transform 1 0 34500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_383
timestamp 1649977179
transform 1 0 36340 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_397
timestamp 1649977179
transform 1 0 37628 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_400
timestamp 1649977179
transform 1 0 37904 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_406
timestamp 1649977179
transform 1 0 38456 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_162
timestamp 1649977179
transform 1 0 16008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_168
timestamp 1649977179
transform 1 0 16560 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_176
timestamp 1649977179
transform 1 0 17296 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_188
timestamp 1649977179
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_201
timestamp 1649977179
transform 1 0 19596 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_207
timestamp 1649977179
transform 1 0 20148 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_214
timestamp 1649977179
transform 1 0 20792 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_222
timestamp 1649977179
transform 1 0 21528 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_241
timestamp 1649977179
transform 1 0 23276 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1649977179
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_291
timestamp 1649977179
transform 1 0 27876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 1649977179
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_347
timestamp 1649977179
transform 1 0 33028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_359
timestamp 1649977179
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_395
timestamp 1649977179
transform 1 0 37444 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_116
timestamp 1649977179
transform 1 0 11776 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_128
timestamp 1649977179
transform 1 0 12880 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_140
timestamp 1649977179
transform 1 0 13984 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_171
timestamp 1649977179
transform 1 0 16836 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_183
timestamp 1649977179
transform 1 0 17940 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_187
timestamp 1649977179
transform 1 0 18308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_201
timestamp 1649977179
transform 1 0 19596 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_209
timestamp 1649977179
transform 1 0 20332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_241
timestamp 1649977179
transform 1 0 23276 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_262
timestamp 1649977179
transform 1 0 25208 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1649977179
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_297
timestamp 1649977179
transform 1 0 28428 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_314
timestamp 1649977179
transform 1 0 29992 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_326
timestamp 1649977179
transform 1 0 31096 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1649977179
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_375
timestamp 1649977179
transform 1 0 35604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_387
timestamp 1649977179
transform 1 0 36708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1649977179
transform 1 0 38180 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1649977179
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_151
timestamp 1649977179
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_157
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_164
timestamp 1649977179
transform 1 0 16192 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_171
timestamp 1649977179
transform 1 0 16836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_178
timestamp 1649977179
transform 1 0 17480 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_185
timestamp 1649977179
transform 1 0 18124 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_200
timestamp 1649977179
transform 1 0 19504 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_212
timestamp 1649977179
transform 1 0 20608 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_240
timestamp 1649977179
transform 1 0 23184 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_261
timestamp 1649977179
transform 1 0 25116 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_278
timestamp 1649977179
transform 1 0 26680 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_290
timestamp 1649977179
transform 1 0 27784 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_302
timestamp 1649977179
transform 1 0 28888 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_317
timestamp 1649977179
transform 1 0 30268 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_334
timestamp 1649977179
transform 1 0 31832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_354
timestamp 1649977179
transform 1 0 33672 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1649977179
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_381
timestamp 1649977179
transform 1 0 36156 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_385
timestamp 1649977179
transform 1 0 36524 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1649977179
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_160
timestamp 1649977179
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_179
timestamp 1649977179
transform 1 0 17572 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_194
timestamp 1649977179
transform 1 0 18952 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_203
timestamp 1649977179
transform 1 0 19780 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_209
timestamp 1649977179
transform 1 0 20332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_241
timestamp 1649977179
transform 1 0 23276 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_266
timestamp 1649977179
transform 1 0 25576 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1649977179
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_298
timestamp 1649977179
transform 1 0 28520 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_310
timestamp 1649977179
transform 1 0 29624 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_322
timestamp 1649977179
transform 1 0 30728 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1649977179
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_354
timestamp 1649977179
transform 1 0 33672 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_366
timestamp 1649977179
transform 1 0 34776 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_378
timestamp 1649977179
transform 1 0 35880 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1649977179
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_151
timestamp 1649977179
transform 1 0 14996 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_166
timestamp 1649977179
transform 1 0 16376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_174
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_181
timestamp 1649977179
transform 1 0 17756 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_188
timestamp 1649977179
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1649977179
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_208
timestamp 1649977179
transform 1 0 20240 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_220
timestamp 1649977179
transform 1 0 21344 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_239
timestamp 1649977179
transform 1 0 23092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_284
timestamp 1649977179
transform 1 0 27232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1649977179
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_327
timestamp 1649977179
transform 1 0 31188 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_339
timestamp 1649977179
transform 1 0 32292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_351
timestamp 1649977179
transform 1 0 33396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_396
timestamp 1649977179
transform 1 0 37536 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_404
timestamp 1649977179
transform 1 0 38272 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_155
timestamp 1649977179
transform 1 0 15364 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_174
timestamp 1649977179
transform 1 0 17112 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_185
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_188
timestamp 1649977179
transform 1 0 18400 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_197
timestamp 1649977179
transform 1 0 19228 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_206
timestamp 1649977179
transform 1 0 20056 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_215
timestamp 1649977179
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_241
timestamp 1649977179
transform 1 0 23276 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_303
timestamp 1649977179
transform 1 0 28980 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_323
timestamp 1649977179
transform 1 0 30820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_353
timestamp 1649977179
transform 1 0 33580 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1649977179
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_396
timestamp 1649977179
transform 1 0 37536 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_404
timestamp 1649977179
transform 1 0 38272 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_147
timestamp 1649977179
transform 1 0 14628 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_155
timestamp 1649977179
transform 1 0 15364 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_158
timestamp 1649977179
transform 1 0 15640 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_164
timestamp 1649977179
transform 1 0 16192 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_173
timestamp 1649977179
transform 1 0 17020 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_179
timestamp 1649977179
transform 1 0 17572 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_185
timestamp 1649977179
transform 1 0 18124 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_200
timestamp 1649977179
transform 1 0 19504 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_207
timestamp 1649977179
transform 1 0 20148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_219
timestamp 1649977179
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_239
timestamp 1649977179
transform 1 0 23092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_270
timestamp 1649977179
transform 1 0 25944 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_290
timestamp 1649977179
transform 1 0 27784 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1649977179
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_343
timestamp 1649977179
transform 1 0 32660 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_355
timestamp 1649977179
transform 1 0 33764 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_385
timestamp 1649977179
transform 1 0 36524 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_403
timestamp 1649977179
transform 1 0 38180 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1649977179
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_172
timestamp 1649977179
transform 1 0 16928 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_183
timestamp 1649977179
transform 1 0 17940 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1649977179
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_192
timestamp 1649977179
transform 1 0 18768 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_204
timestamp 1649977179
transform 1 0 19872 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_210
timestamp 1649977179
transform 1 0 20424 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1649977179
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_266
timestamp 1649977179
transform 1 0 25576 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1649977179
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_381
timestamp 1649977179
transform 1 0 36156 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_159
timestamp 1649977179
transform 1 0 15732 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_167
timestamp 1649977179
transform 1 0 16468 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 1649977179
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_199
timestamp 1649977179
transform 1 0 19412 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_207
timestamp 1649977179
transform 1 0 20148 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_212
timestamp 1649977179
transform 1 0 20608 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_218
timestamp 1649977179
transform 1 0 21160 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_230
timestamp 1649977179
transform 1 0 22264 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_236
timestamp 1649977179
transform 1 0 22816 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1649977179
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_264
timestamp 1649977179
transform 1 0 25392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_270
timestamp 1649977179
transform 1 0 25944 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_276
timestamp 1649977179
transform 1 0 26496 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_288
timestamp 1649977179
transform 1 0 27600 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_296
timestamp 1649977179
transform 1 0 28336 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_336
timestamp 1649977179
transform 1 0 32016 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_352
timestamp 1649977179
transform 1 0 33488 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_373
timestamp 1649977179
transform 1 0 35420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_390
timestamp 1649977179
transform 1 0 36984 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_402
timestamp 1649977179
transform 1 0 38088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_406
timestamp 1649977179
transform 1 0 38456 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1649977179
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_176
timestamp 1649977179
transform 1 0 17296 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_182
timestamp 1649977179
transform 1 0 17848 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_188
timestamp 1649977179
transform 1 0 18400 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_196
timestamp 1649977179
transform 1 0 19136 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_208
timestamp 1649977179
transform 1 0 20240 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_216
timestamp 1649977179
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_234
timestamp 1649977179
transform 1 0 22632 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_242
timestamp 1649977179
transform 1 0 23368 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_248
timestamp 1649977179
transform 1 0 23920 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_263
timestamp 1649977179
transform 1 0 25300 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1649977179
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_320
timestamp 1649977179
transform 1 0 30544 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_328
timestamp 1649977179
transform 1 0 31280 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1649977179
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_342
timestamp 1649977179
transform 1 0 32568 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_354
timestamp 1649977179
transform 1 0 33672 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_366
timestamp 1649977179
transform 1 0 34776 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_378
timestamp 1649977179
transform 1 0 35880 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1649977179
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_176
timestamp 1649977179
transform 1 0 17296 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_187
timestamp 1649977179
transform 1 0 18308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_214
timestamp 1649977179
transform 1 0 20792 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_220
timestamp 1649977179
transform 1 0 21344 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_227
timestamp 1649977179
transform 1 0 21988 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_236
timestamp 1649977179
transform 1 0 22816 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1649977179
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_256
timestamp 1649977179
transform 1 0 24656 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_262
timestamp 1649977179
transform 1 0 25208 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_278
timestamp 1649977179
transform 1 0 26680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1649977179
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_381
timestamp 1649977179
transform 1 0 36156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_394
timestamp 1649977179
transform 1 0 37352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_175
timestamp 1649977179
transform 1 0 17204 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_178
timestamp 1649977179
transform 1 0 17480 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_190
timestamp 1649977179
transform 1 0 18584 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_201
timestamp 1649977179
transform 1 0 19596 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_207
timestamp 1649977179
transform 1 0 20148 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1649977179
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_230
timestamp 1649977179
transform 1 0 22264 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_234
timestamp 1649977179
transform 1 0 22632 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_244
timestamp 1649977179
transform 1 0 23552 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_250
timestamp 1649977179
transform 1 0 24104 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_256
timestamp 1649977179
transform 1 0 24656 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_268
timestamp 1649977179
transform 1 0 25760 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1649977179
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_203
timestamp 1649977179
transform 1 0 19780 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_220
timestamp 1649977179
transform 1 0 21344 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_226
timestamp 1649977179
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_232
timestamp 1649977179
transform 1 0 22448 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_244
timestamp 1649977179
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_196
timestamp 1649977179
transform 1 0 19136 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_202
timestamp 1649977179
transform 1 0 19688 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_214
timestamp 1649977179
transform 1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1649977179
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_270
timestamp 1649977179
transform 1 0 25944 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1649977179
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_283
timestamp 1649977179
transform 1 0 27140 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_295
timestamp 1649977179
transform 1 0 28244 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_307
timestamp 1649977179
transform 1 0 29348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_319
timestamp 1649977179
transform 1 0 30452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_331
timestamp 1649977179
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_183
timestamp 1649977179
transform 1 0 17940 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_186
timestamp 1649977179
transform 1 0 18216 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1649977179
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_367
timestamp 1649977179
transform 1 0 34868 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_379
timestamp 1649977179
transform 1 0 35972 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_391
timestamp 1649977179
transform 1 0 37076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_403
timestamp 1649977179
transform 1 0 38180 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_184
timestamp 1649977179
transform 1 0 18032 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_190
timestamp 1649977179
transform 1 0 18584 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_202
timestamp 1649977179
transform 1 0 19688 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_214
timestamp 1649977179
transform 1 0 20792 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1649977179
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_345
timestamp 1649977179
transform 1 0 32844 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_348
timestamp 1649977179
transform 1 0 33120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_368
timestamp 1649977179
transform 1 0 34960 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_380
timestamp 1649977179
transform 1 0 36064 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_239
timestamp 1649977179
transform 1 0 23092 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_385
timestamp 1649977179
transform 1 0 36524 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_397
timestamp 1649977179
transform 1 0 37628 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_405
timestamp 1649977179
transform 1 0 38364 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_213
timestamp 1649977179
transform 1 0 20700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1649977179
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_227
timestamp 1649977179
transform 1 0 21988 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_239
timestamp 1649977179
transform 1 0 23092 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_251
timestamp 1649977179
transform 1 0 24196 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_263
timestamp 1649977179
transform 1 0 25300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 1649977179
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_309
timestamp 1649977179
transform 1 0 29532 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_318
timestamp 1649977179
transform 1 0 30360 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_330
timestamp 1649977179
transform 1 0 31464 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_361
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_367
timestamp 1649977179
transform 1 0 34868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_370
timestamp 1649977179
transform 1 0 35144 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_383
timestamp 1649977179
transform 1 0 36340 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_212
timestamp 1649977179
transform 1 0 20608 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_225
timestamp 1649977179
transform 1 0 21804 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_231
timestamp 1649977179
transform 1 0 22356 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_237
timestamp 1649977179
transform 1 0 22908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1649977179
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1649977179
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_314
timestamp 1649977179
transform 1 0 29992 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_320
timestamp 1649977179
transform 1 0 30544 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_332
timestamp 1649977179
transform 1 0 31648 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_344
timestamp 1649977179
transform 1 0 32752 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_356
timestamp 1649977179
transform 1 0 33856 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_373
timestamp 1649977179
transform 1 0 35420 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_376
timestamp 1649977179
transform 1 0 35696 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1649977179
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_215
timestamp 1649977179
transform 1 0 20884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_227
timestamp 1649977179
transform 1 0 21988 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_239
timestamp 1649977179
transform 1 0 23092 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_251
timestamp 1649977179
transform 1 0 24196 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_263
timestamp 1649977179
transform 1 0 25300 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1649977179
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_297
timestamp 1649977179
transform 1 0 28428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_303
timestamp 1649977179
transform 1 0 28980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_318
timestamp 1649977179
transform 1 0 30360 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_324
timestamp 1649977179
transform 1 0 30912 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_330
timestamp 1649977179
transform 1 0 31464 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1649977179
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_217
timestamp 1649977179
transform 1 0 21068 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_229
timestamp 1649977179
transform 1 0 22172 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_241
timestamp 1649977179
transform 1 0 23276 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1649977179
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_285
timestamp 1649977179
transform 1 0 27324 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_291
timestamp 1649977179
transform 1 0 27876 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_320
timestamp 1649977179
transform 1 0 30544 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_339
timestamp 1649977179
transform 1 0 32292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_351
timestamp 1649977179
transform 1 0 33396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_369
timestamp 1649977179
transform 1 0 35052 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_372
timestamp 1649977179
transform 1 0 35328 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_385
timestamp 1649977179
transform 1 0 36524 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_391
timestamp 1649977179
transform 1 0 37076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_403
timestamp 1649977179
transform 1 0 38180 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1649977179
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_283
timestamp 1649977179
transform 1 0 27140 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_300
timestamp 1649977179
transform 1 0 28704 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_306
timestamp 1649977179
transform 1 0 29256 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_312
timestamp 1649977179
transform 1 0 29808 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_318
timestamp 1649977179
transform 1 0 30360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_322
timestamp 1649977179
transform 1 0 30728 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1649977179
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_339
timestamp 1649977179
transform 1 0 32292 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_345
timestamp 1649977179
transform 1 0 32844 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_357
timestamp 1649977179
transform 1 0 33948 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_362
timestamp 1649977179
transform 1 0 34408 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_376
timestamp 1649977179
transform 1 0 35696 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_230
timestamp 1649977179
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_236
timestamp 1649977179
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_242
timestamp 1649977179
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1649977179
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_268
timestamp 1649977179
transform 1 0 25760 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_281
timestamp 1649977179
transform 1 0 26956 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_287
timestamp 1649977179
transform 1 0 27508 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_293
timestamp 1649977179
transform 1 0 28060 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_302
timestamp 1649977179
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_317
timestamp 1649977179
transform 1 0 30268 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_329
timestamp 1649977179
transform 1 0 31372 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_341
timestamp 1649977179
transform 1 0 32476 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_349
timestamp 1649977179
transform 1 0 33212 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1649977179
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_374
timestamp 1649977179
transform 1 0 35512 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_387
timestamp 1649977179
transform 1 0 36708 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_393
timestamp 1649977179
transform 1 0 37260 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1649977179
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_213
timestamp 1649977179
transform 1 0 20700 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1649977179
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_234
timestamp 1649977179
transform 1 0 22632 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_243
timestamp 1649977179
transform 1 0 23460 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_255
timestamp 1649977179
transform 1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_263
timestamp 1649977179
transform 1 0 25300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1649977179
transform 1 0 25852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1649977179
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_285
timestamp 1649977179
transform 1 0 27324 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_292
timestamp 1649977179
transform 1 0 27968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_299
timestamp 1649977179
transform 1 0 28612 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_307
timestamp 1649977179
transform 1 0 29348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_315
timestamp 1649977179
transform 1 0 30084 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_323
timestamp 1649977179
transform 1 0 30820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_340
timestamp 1649977179
transform 1 0 32384 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_348
timestamp 1649977179
transform 1 0 33120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_352
timestamp 1649977179
transform 1 0 33488 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_367
timestamp 1649977179
transform 1 0 34868 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_380
timestamp 1649977179
transform 1 0 36064 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_180
timestamp 1649977179
transform 1 0 17664 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1649977179
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_205
timestamp 1649977179
transform 1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_218
timestamp 1649977179
transform 1 0 21160 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_222
timestamp 1649977179
transform 1 0 21528 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_225
timestamp 1649977179
transform 1 0 21804 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_231
timestamp 1649977179
transform 1 0 22356 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_241
timestamp 1649977179
transform 1 0 23276 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_247
timestamp 1649977179
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_258
timestamp 1649977179
transform 1 0 24840 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_279
timestamp 1649977179
transform 1 0 26772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_291
timestamp 1649977179
transform 1 0 27876 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_298
timestamp 1649977179
transform 1 0 28520 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1649977179
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_311
timestamp 1649977179
transform 1 0 29716 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_317
timestamp 1649977179
transform 1 0 30268 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_327
timestamp 1649977179
transform 1 0 31188 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_334
timestamp 1649977179
transform 1 0 31832 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_342
timestamp 1649977179
transform 1 0 32568 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_351
timestamp 1649977179
transform 1 0 33396 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_355
timestamp 1649977179
transform 1 0 33764 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_358
timestamp 1649977179
transform 1 0 34040 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_370
timestamp 1649977179
transform 1 0 35144 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_379
timestamp 1649977179
transform 1 0 35972 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_387
timestamp 1649977179
transform 1 0 36708 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_391
timestamp 1649977179
transform 1 0 37076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_403
timestamp 1649977179
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1649977179
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_178
timestamp 1649977179
transform 1 0 17480 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_184
timestamp 1649977179
transform 1 0 18032 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_190
timestamp 1649977179
transform 1 0 18584 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_194
timestamp 1649977179
transform 1 0 18952 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_200
timestamp 1649977179
transform 1 0 19504 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_210
timestamp 1649977179
transform 1 0 20424 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1649977179
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_238
timestamp 1649977179
transform 1 0 23000 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_247
timestamp 1649977179
transform 1 0 23828 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_258
timestamp 1649977179
transform 1 0 24840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1649977179
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_283
timestamp 1649977179
transform 1 0 27140 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_289
timestamp 1649977179
transform 1 0 27692 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_292
timestamp 1649977179
transform 1 0 27968 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_309
timestamp 1649977179
transform 1 0 29532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_315
timestamp 1649977179
transform 1 0 30084 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_328
timestamp 1649977179
transform 1 0 31280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_346
timestamp 1649977179
transform 1 0 32936 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_352
timestamp 1649977179
transform 1 0 33488 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_367
timestamp 1649977179
transform 1 0 34868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_379
timestamp 1649977179
transform 1 0 35972 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_126
timestamp 1649977179
transform 1 0 12696 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1649977179
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_145
timestamp 1649977179
transform 1 0 14444 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_156
timestamp 1649977179
transform 1 0 15456 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_168
timestamp 1649977179
transform 1 0 16560 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_174
timestamp 1649977179
transform 1 0 17112 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_183
timestamp 1649977179
transform 1 0 17940 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1649977179
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_206
timestamp 1649977179
transform 1 0 20056 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_212
timestamp 1649977179
transform 1 0 20608 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_219
timestamp 1649977179
transform 1 0 21252 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_227
timestamp 1649977179
transform 1 0 21988 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_237
timestamp 1649977179
transform 1 0 22908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_243
timestamp 1649977179
transform 1 0 23460 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_255
timestamp 1649977179
transform 1 0 24564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_261
timestamp 1649977179
transform 1 0 25116 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_267
timestamp 1649977179
transform 1 0 25668 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_279
timestamp 1649977179
transform 1 0 26772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_294
timestamp 1649977179
transform 1 0 28152 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_298
timestamp 1649977179
transform 1 0 28520 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_302
timestamp 1649977179
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_314
timestamp 1649977179
transform 1 0 29992 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_328
timestamp 1649977179
transform 1 0 31280 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_332
timestamp 1649977179
transform 1 0 31648 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_338
timestamp 1649977179
transform 1 0 32200 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_353
timestamp 1649977179
transform 1 0 33580 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_359
timestamp 1649977179
transform 1 0 34132 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_370
timestamp 1649977179
transform 1 0 35144 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_386
timestamp 1649977179
transform 1 0 36616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_392
timestamp 1649977179
transform 1 0 37168 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_403
timestamp 1649977179
transform 1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1649977179
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1649977179
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1649977179
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_96
timestamp 1649977179
transform 1 0 9936 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1649977179
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_122
timestamp 1649977179
transform 1 0 12328 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_128
timestamp 1649977179
transform 1 0 12880 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_141
timestamp 1649977179
transform 1 0 14076 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_154
timestamp 1649977179
transform 1 0 15272 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_160
timestamp 1649977179
transform 1 0 15824 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_171
timestamp 1649977179
transform 1 0 16836 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_184
timestamp 1649977179
transform 1 0 18032 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_190
timestamp 1649977179
transform 1 0 18584 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_198
timestamp 1649977179
transform 1 0 19320 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_215
timestamp 1649977179
transform 1 0 20884 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_234
timestamp 1649977179
transform 1 0 22632 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_238
timestamp 1649977179
transform 1 0 23000 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_242
timestamp 1649977179
transform 1 0 23368 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_248
timestamp 1649977179
transform 1 0 23920 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_254
timestamp 1649977179
transform 1 0 24472 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_266
timestamp 1649977179
transform 1 0 25576 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1649977179
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_305
timestamp 1649977179
transform 1 0 29164 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_312
timestamp 1649977179
transform 1 0 29808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_318
timestamp 1649977179
transform 1 0 30360 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_326
timestamp 1649977179
transform 1 0 31096 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1649977179
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_339
timestamp 1649977179
transform 1 0 32292 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_350
timestamp 1649977179
transform 1 0 33304 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_356
timestamp 1649977179
transform 1 0 33856 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_362
timestamp 1649977179
transform 1 0 34408 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_382
timestamp 1649977179
transform 1 0 36248 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_388
timestamp 1649977179
transform 1 0 36800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_403
timestamp 1649977179
transform 1 0 38180 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_94
timestamp 1649977179
transform 1 0 9752 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_100
timestamp 1649977179
transform 1 0 10304 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_106
timestamp 1649977179
transform 1 0 10856 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_123
timestamp 1649977179
transform 1 0 12420 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_129
timestamp 1649977179
transform 1 0 12972 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_135
timestamp 1649977179
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_143
timestamp 1649977179
transform 1 0 14260 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_151
timestamp 1649977179
transform 1 0 14996 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_161
timestamp 1649977179
transform 1 0 15916 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_169
timestamp 1649977179
transform 1 0 16652 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_179
timestamp 1649977179
transform 1 0 17572 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1649977179
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_201
timestamp 1649977179
transform 1 0 19596 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_207
timestamp 1649977179
transform 1 0 20148 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_213
timestamp 1649977179
transform 1 0 20700 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_219
timestamp 1649977179
transform 1 0 21252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_223
timestamp 1649977179
transform 1 0 21620 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_226
timestamp 1649977179
transform 1 0 21896 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_235
timestamp 1649977179
transform 1 0 22724 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_241
timestamp 1649977179
transform 1 0 23276 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_247
timestamp 1649977179
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_269
timestamp 1649977179
transform 1 0 25852 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_325
timestamp 1649977179
transform 1 0 31004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_353
timestamp 1649977179
transform 1 0 33580 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_368
timestamp 1649977179
transform 1 0 34960 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_383
timestamp 1649977179
transform 1 0 36340 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_403
timestamp 1649977179
transform 1 0 38180 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_90
timestamp 1649977179
transform 1 0 9384 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_100
timestamp 1649977179
transform 1 0 10304 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_106
timestamp 1649977179
transform 1 0 10856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_121
timestamp 1649977179
transform 1 0 12236 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_155
timestamp 1649977179
transform 1 0 15364 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_158
timestamp 1649977179
transform 1 0 15640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1649977179
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_178
timestamp 1649977179
transform 1 0 17480 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_188
timestamp 1649977179
transform 1 0 18400 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_194
timestamp 1649977179
transform 1 0 18952 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_202
timestamp 1649977179
transform 1 0 19688 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_215
timestamp 1649977179
transform 1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_232
timestamp 1649977179
transform 1 0 22448 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_244
timestamp 1649977179
transform 1 0 23552 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_266
timestamp 1649977179
transform 1 0 25576 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1649977179
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_319
timestamp 1649977179
transform 1 0 30452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_331
timestamp 1649977179
transform 1 0 31556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_353
timestamp 1649977179
transform 1 0 33580 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_365
timestamp 1649977179
transform 1 0 34684 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_371
timestamp 1649977179
transform 1 0 35236 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_388
timestamp 1649977179
transform 1 0 36800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_402
timestamp 1649977179
transform 1 0 38088 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_406
timestamp 1649977179
transform 1 0 38456 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_96
timestamp 1649977179
transform 1 0 9936 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_102
timestamp 1649977179
transform 1 0 10488 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_111
timestamp 1649977179
transform 1 0 11316 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_118
timestamp 1649977179
transform 1 0 11960 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_130
timestamp 1649977179
transform 1 0 13064 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_147
timestamp 1649977179
transform 1 0 14628 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_151
timestamp 1649977179
transform 1 0 14996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_163
timestamp 1649977179
transform 1 0 16100 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_166
timestamp 1649977179
transform 1 0 16376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_175
timestamp 1649977179
transform 1 0 17204 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_181
timestamp 1649977179
transform 1 0 17756 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_191
timestamp 1649977179
transform 1 0 18676 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_206
timestamp 1649977179
transform 1 0 20056 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_212
timestamp 1649977179
transform 1 0 20608 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_227
timestamp 1649977179
transform 1 0 21988 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_239
timestamp 1649977179
transform 1 0 23092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_291
timestamp 1649977179
transform 1 0 27876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_303
timestamp 1649977179
transform 1 0 28980 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_347
timestamp 1649977179
transform 1 0 33028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_359
timestamp 1649977179
transform 1 0 34132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_371
timestamp 1649977179
transform 1 0 35236 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_375
timestamp 1649977179
transform 1 0 35604 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_403
timestamp 1649977179
transform 1 0 38180 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_77
timestamp 1649977179
transform 1 0 8188 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_84
timestamp 1649977179
transform 1 0 8832 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_100
timestamp 1649977179
transform 1 0 10304 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_117
timestamp 1649977179
transform 1 0 11868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_121
timestamp 1649977179
transform 1 0 12236 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_131
timestamp 1649977179
transform 1 0 13156 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_143
timestamp 1649977179
transform 1 0 14260 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_153
timestamp 1649977179
transform 1 0 15180 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_156
timestamp 1649977179
transform 1 0 15456 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1649977179
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_173
timestamp 1649977179
transform 1 0 17020 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_182
timestamp 1649977179
transform 1 0 17848 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_186
timestamp 1649977179
transform 1 0 18216 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_189
timestamp 1649977179
transform 1 0 18492 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_198
timestamp 1649977179
transform 1 0 19320 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_209
timestamp 1649977179
transform 1 0 20332 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_215
timestamp 1649977179
transform 1 0 20884 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_231
timestamp 1649977179
transform 1 0 22356 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_269
timestamp 1649977179
transform 1 0 25852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1649977179
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_297
timestamp 1649977179
transform 1 0 28428 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_309
timestamp 1649977179
transform 1 0 29532 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_328
timestamp 1649977179
transform 1 0 31280 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_353
timestamp 1649977179
transform 1 0 33580 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_105
timestamp 1649977179
transform 1 0 10764 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_111
timestamp 1649977179
transform 1 0 11316 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_117
timestamp 1649977179
transform 1 0 11868 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_127
timestamp 1649977179
transform 1 0 12788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_150
timestamp 1649977179
transform 1 0 14904 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_159
timestamp 1649977179
transform 1 0 15732 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_168
timestamp 1649977179
transform 1 0 16560 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_180
timestamp 1649977179
transform 1 0 17664 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_185
timestamp 1649977179
transform 1 0 18124 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1649977179
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_199
timestamp 1649977179
transform 1 0 19412 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_205
timestamp 1649977179
transform 1 0 19964 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_214
timestamp 1649977179
transform 1 0 20792 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_222
timestamp 1649977179
transform 1 0 21528 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_226
timestamp 1649977179
transform 1 0 21896 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_269
timestamp 1649977179
transform 1 0 25852 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_290
timestamp 1649977179
transform 1 0 27784 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_302
timestamp 1649977179
transform 1 0 28888 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_341
timestamp 1649977179
transform 1 0 32476 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1649977179
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_373
timestamp 1649977179
transform 1 0 35420 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_391
timestamp 1649977179
transform 1 0 37076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_403
timestamp 1649977179
transform 1 0 38180 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_89
timestamp 1649977179
transform 1 0 9292 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_97
timestamp 1649977179
transform 1 0 10028 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_106
timestamp 1649977179
transform 1 0 10856 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_122
timestamp 1649977179
transform 1 0 12328 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_131
timestamp 1649977179
transform 1 0 13156 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_151
timestamp 1649977179
transform 1 0 14996 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1649977179
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_172
timestamp 1649977179
transform 1 0 16928 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_184
timestamp 1649977179
transform 1 0 18032 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_197
timestamp 1649977179
transform 1 0 19228 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_205
timestamp 1649977179
transform 1 0 19964 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_209
timestamp 1649977179
transform 1 0 20332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1649977179
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_265
timestamp 1649977179
transform 1 0 25484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_277
timestamp 1649977179
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_315
timestamp 1649977179
transform 1 0 30084 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_327
timestamp 1649977179
transform 1 0 31188 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1649977179
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_357
timestamp 1649977179
transform 1 0 33948 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_374
timestamp 1649977179
transform 1 0 35512 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_386
timestamp 1649977179
transform 1 0 36616 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_95
timestamp 1649977179
transform 1 0 9844 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_108
timestamp 1649977179
transform 1 0 11040 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_117
timestamp 1649977179
transform 1 0 11868 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_123
timestamp 1649977179
transform 1 0 12420 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_129
timestamp 1649977179
transform 1 0 12972 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_137
timestamp 1649977179
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_146
timestamp 1649977179
transform 1 0 14536 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_154
timestamp 1649977179
transform 1 0 15272 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_160
timestamp 1649977179
transform 1 0 15824 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_166
timestamp 1649977179
transform 1 0 16376 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_172
timestamp 1649977179
transform 1 0 16928 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_178
timestamp 1649977179
transform 1 0 17480 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_190
timestamp 1649977179
transform 1 0 18584 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_217
timestamp 1649977179
transform 1 0 21068 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_221
timestamp 1649977179
transform 1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_227
timestamp 1649977179
transform 1 0 21988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_239
timestamp 1649977179
transform 1 0 23092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_259
timestamp 1649977179
transform 1 0 24932 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_276
timestamp 1649977179
transform 1 0 26496 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1649977179
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_340
timestamp 1649977179
transform 1 0 32384 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_352
timestamp 1649977179
transform 1 0 33488 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_385
timestamp 1649977179
transform 1 0 36524 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_403
timestamp 1649977179
transform 1 0 38180 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1649977179
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_95
timestamp 1649977179
transform 1 0 9844 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_101
timestamp 1649977179
transform 1 0 10396 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_107
timestamp 1649977179
transform 1 0 10948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_115
timestamp 1649977179
transform 1 0 11684 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_119
timestamp 1649977179
transform 1 0 12052 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_123
timestamp 1649977179
transform 1 0 12420 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_132
timestamp 1649977179
transform 1 0 13248 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_144
timestamp 1649977179
transform 1 0 14352 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_152
timestamp 1649977179
transform 1 0 15088 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_158
timestamp 1649977179
transform 1 0 15640 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1649977179
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_193
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_199
timestamp 1649977179
transform 1 0 19412 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_203
timestamp 1649977179
transform 1 0 19780 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1649977179
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_230
timestamp 1649977179
transform 1 0 22264 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_236
timestamp 1649977179
transform 1 0 22816 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_248
timestamp 1649977179
transform 1 0 23920 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_252
timestamp 1649977179
transform 1 0 24288 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_269
timestamp 1649977179
transform 1 0 25852 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 1649977179
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_289
timestamp 1649977179
transform 1 0 27692 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_308
timestamp 1649977179
transform 1 0 29440 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_320
timestamp 1649977179
transform 1 0 30544 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1649977179
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1649977179
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1649977179
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_130
timestamp 1649977179
transform 1 0 13064 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1649977179
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_144
timestamp 1649977179
transform 1 0 14352 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_152
timestamp 1649977179
transform 1 0 15088 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_162
timestamp 1649977179
transform 1 0 16008 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_168
timestamp 1649977179
transform 1 0 16560 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_172
timestamp 1649977179
transform 1 0 16928 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_176
timestamp 1649977179
transform 1 0 17296 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_188
timestamp 1649977179
transform 1 0 18400 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_229
timestamp 1649977179
transform 1 0 22172 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_236
timestamp 1649977179
transform 1 0 22816 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_242
timestamp 1649977179
transform 1 0 23368 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1649977179
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_269
timestamp 1649977179
transform 1 0 25852 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_281
timestamp 1649977179
transform 1 0 26956 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_293
timestamp 1649977179
transform 1 0 28060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_305
timestamp 1649977179
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_337
timestamp 1649977179
transform 1 0 32108 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_349
timestamp 1649977179
transform 1 0 33212 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_361
timestamp 1649977179
transform 1 0 34316 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_383
timestamp 1649977179
transform 1 0 36340 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_403
timestamp 1649977179
transform 1 0 38180 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1649977179
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_118
timestamp 1649977179
transform 1 0 11960 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_132
timestamp 1649977179
transform 1 0 13248 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_138
timestamp 1649977179
transform 1 0 13800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_146
timestamp 1649977179
transform 1 0 14536 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_157
timestamp 1649977179
transform 1 0 15548 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1649977179
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_177
timestamp 1649977179
transform 1 0 17388 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_187
timestamp 1649977179
transform 1 0 18308 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_199
timestamp 1649977179
transform 1 0 19412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_211
timestamp 1649977179
transform 1 0 20516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_227
timestamp 1649977179
transform 1 0 21988 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_233
timestamp 1649977179
transform 1 0 22540 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_245
timestamp 1649977179
transform 1 0 23644 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_269
timestamp 1649977179
transform 1 0 25852 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1649977179
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_298
timestamp 1649977179
transform 1 0 28520 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_318
timestamp 1649977179
transform 1 0 30360 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_330
timestamp 1649977179
transform 1 0 31464 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_368
timestamp 1649977179
transform 1 0 34960 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_380
timestamp 1649977179
transform 1 0 36064 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1649977179
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_115
timestamp 1649977179
transform 1 0 11684 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_128
timestamp 1649977179
transform 1 0 12880 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_180
timestamp 1649977179
transform 1 0 17664 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_207
timestamp 1649977179
transform 1 0 20148 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_216
timestamp 1649977179
transform 1 0 20976 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_228
timestamp 1649977179
transform 1 0 22080 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_240
timestamp 1649977179
transform 1 0 23184 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_291
timestamp 1649977179
transform 1 0 27876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1649977179
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_340
timestamp 1649977179
transform 1 0 32384 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_352
timestamp 1649977179
transform 1 0 33488 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_385
timestamp 1649977179
transform 1 0 36524 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_397
timestamp 1649977179
transform 1 0 37628 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_405
timestamp 1649977179
transform 1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1649977179
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_172
timestamp 1649977179
transform 1 0 16928 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_180
timestamp 1649977179
transform 1 0 17664 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_184
timestamp 1649977179
transform 1 0 18032 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_188
timestamp 1649977179
transform 1 0 18400 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_196
timestamp 1649977179
transform 1 0 19136 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_208
timestamp 1649977179
transform 1 0 20240 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_213
timestamp 1649977179
transform 1 0 20700 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_221
timestamp 1649977179
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_234
timestamp 1649977179
transform 1 0 22632 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_240
timestamp 1649977179
transform 1 0 23184 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_268
timestamp 1649977179
transform 1 0 25760 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_297
timestamp 1649977179
transform 1 0 28428 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_303
timestamp 1649977179
transform 1 0 28980 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_320
timestamp 1649977179
transform 1 0 30544 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1649977179
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_381
timestamp 1649977179
transform 1 0 36156 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_389
timestamp 1649977179
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_136
timestamp 1649977179
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_147
timestamp 1649977179
transform 1 0 14628 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_155
timestamp 1649977179
transform 1 0 15364 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_165
timestamp 1649977179
transform 1 0 16284 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_172
timestamp 1649977179
transform 1 0 16928 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_184
timestamp 1649977179
transform 1 0 18032 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_199
timestamp 1649977179
transform 1 0 19412 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_211
timestamp 1649977179
transform 1 0 20516 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_223
timestamp 1649977179
transform 1 0 21620 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_230
timestamp 1649977179
transform 1 0 22264 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_236
timestamp 1649977179
transform 1 0 22816 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_240
timestamp 1649977179
transform 1 0 23184 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_269
timestamp 1649977179
transform 1 0 25852 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_281
timestamp 1649977179
transform 1 0 26956 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_293
timestamp 1649977179
transform 1 0 28060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_305
timestamp 1649977179
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_311
timestamp 1649977179
transform 1 0 29716 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_319
timestamp 1649977179
transform 1 0 30452 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_324
timestamp 1649977179
transform 1 0 30912 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_344
timestamp 1649977179
transform 1 0 32752 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_356
timestamp 1649977179
transform 1 0 33856 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_367
timestamp 1649977179
transform 1 0 34868 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_373
timestamp 1649977179
transform 1 0 35420 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_385
timestamp 1649977179
transform 1 0 36524 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_403
timestamp 1649977179
transform 1 0 38180 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1649977179
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_55_124
timestamp 1649977179
transform 1 0 12512 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_130
timestamp 1649977179
transform 1 0 13064 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_135
timestamp 1649977179
transform 1 0 13524 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_145
timestamp 1649977179
transform 1 0 14444 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_151
timestamp 1649977179
transform 1 0 14996 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_163
timestamp 1649977179
transform 1 0 16100 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_185
timestamp 1649977179
transform 1 0 18124 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_188
timestamp 1649977179
transform 1 0 18400 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_197
timestamp 1649977179
transform 1 0 19228 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_201
timestamp 1649977179
transform 1 0 19596 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_227
timestamp 1649977179
transform 1 0 21988 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_233
timestamp 1649977179
transform 1 0 22540 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_255
timestamp 1649977179
transform 1 0 24564 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_272
timestamp 1649977179
transform 1 0 26128 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_289
timestamp 1649977179
transform 1 0 27692 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_306
timestamp 1649977179
transform 1 0 29256 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_326
timestamp 1649977179
transform 1 0 31096 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1649977179
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_367
timestamp 1649977179
transform 1 0 34868 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_384
timestamp 1649977179
transform 1 0 36432 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_93
timestamp 1649977179
transform 1 0 9660 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_96
timestamp 1649977179
transform 1 0 9936 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_108
timestamp 1649977179
transform 1 0 11040 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_120
timestamp 1649977179
transform 1 0 12144 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_124
timestamp 1649977179
transform 1 0 12512 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_128
timestamp 1649977179
transform 1 0 12880 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_134
timestamp 1649977179
transform 1 0 13432 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_143
timestamp 1649977179
transform 1 0 14260 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_155
timestamp 1649977179
transform 1 0 15364 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_167
timestamp 1649977179
transform 1 0 16468 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_179
timestamp 1649977179
transform 1 0 17572 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_199
timestamp 1649977179
transform 1 0 19412 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_211
timestamp 1649977179
transform 1 0 20516 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_223
timestamp 1649977179
transform 1 0 21620 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_231
timestamp 1649977179
transform 1 0 22356 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_236
timestamp 1649977179
transform 1 0 22816 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_242
timestamp 1649977179
transform 1 0 23368 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1649977179
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_269
timestamp 1649977179
transform 1 0 25852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_296
timestamp 1649977179
transform 1 0 28336 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_317
timestamp 1649977179
transform 1 0 30268 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_335
timestamp 1649977179
transform 1 0 31924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_355
timestamp 1649977179
transform 1 0 33764 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_85
timestamp 1649977179
transform 1 0 8924 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_92
timestamp 1649977179
transform 1 0 9568 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_100
timestamp 1649977179
transform 1 0 10304 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_106
timestamp 1649977179
transform 1 0 10856 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_115
timestamp 1649977179
transform 1 0 11684 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_123
timestamp 1649977179
transform 1 0 12420 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_130
timestamp 1649977179
transform 1 0 13064 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_138
timestamp 1649977179
transform 1 0 13800 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_143
timestamp 1649977179
transform 1 0 14260 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_151
timestamp 1649977179
transform 1 0 14996 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_163
timestamp 1649977179
transform 1 0 16100 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_172
timestamp 1649977179
transform 1 0 16928 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_57_180
timestamp 1649977179
transform 1 0 17664 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_189
timestamp 1649977179
transform 1 0 18492 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_201
timestamp 1649977179
transform 1 0 19596 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_211
timestamp 1649977179
transform 1 0 20516 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_234
timestamp 1649977179
transform 1 0 22632 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_247
timestamp 1649977179
transform 1 0 23828 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_253
timestamp 1649977179
transform 1 0 24380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_265
timestamp 1649977179
transform 1 0 25484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_277
timestamp 1649977179
transform 1 0 26588 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_319
timestamp 1649977179
transform 1 0 30452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_331
timestamp 1649977179
transform 1 0 31556 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_375
timestamp 1649977179
transform 1 0 35604 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_379
timestamp 1649977179
transform 1 0 35972 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_383
timestamp 1649977179
transform 1 0 36340 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_91
timestamp 1649977179
transform 1 0 9476 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_104
timestamp 1649977179
transform 1 0 10672 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_112
timestamp 1649977179
transform 1 0 11408 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_123
timestamp 1649977179
transform 1 0 12420 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_132
timestamp 1649977179
transform 1 0 13248 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_58_145
timestamp 1649977179
transform 1 0 14444 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_156
timestamp 1649977179
transform 1 0 15456 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_164
timestamp 1649977179
transform 1 0 16192 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_171
timestamp 1649977179
transform 1 0 16836 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_179
timestamp 1649977179
transform 1 0 17572 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_188
timestamp 1649977179
transform 1 0 18400 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_199
timestamp 1649977179
transform 1 0 19412 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_211
timestamp 1649977179
transform 1 0 20516 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_216
timestamp 1649977179
transform 1 0 20976 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_223
timestamp 1649977179
transform 1 0 21620 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_230
timestamp 1649977179
transform 1 0 22264 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_236
timestamp 1649977179
transform 1 0 22816 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_246
timestamp 1649977179
transform 1 0 23736 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_255
timestamp 1649977179
transform 1 0 24564 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_261
timestamp 1649977179
transform 1 0 25116 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_267
timestamp 1649977179
transform 1 0 25668 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_273
timestamp 1649977179
transform 1 0 26220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_294
timestamp 1649977179
transform 1 0 28152 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1649977179
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_347
timestamp 1649977179
transform 1 0 33028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_359
timestamp 1649977179
transform 1 0 34132 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_381
timestamp 1649977179
transform 1 0 36156 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_403
timestamp 1649977179
transform 1 0 38180 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1649977179
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1649977179
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1649977179
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_89
timestamp 1649977179
transform 1 0 9292 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_101
timestamp 1649977179
transform 1 0 10396 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_107
timestamp 1649977179
transform 1 0 10948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_117
timestamp 1649977179
transform 1 0 11868 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_122
timestamp 1649977179
transform 1 0 12328 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_131
timestamp 1649977179
transform 1 0 13156 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_138
timestamp 1649977179
transform 1 0 13800 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_151
timestamp 1649977179
transform 1 0 14996 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_157
timestamp 1649977179
transform 1 0 15548 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_160
timestamp 1649977179
transform 1 0 15824 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_203
timestamp 1649977179
transform 1 0 19780 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_207
timestamp 1649977179
transform 1 0 20148 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_228
timestamp 1649977179
transform 1 0 22080 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_232
timestamp 1649977179
transform 1 0 22448 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_236
timestamp 1649977179
transform 1 0 22816 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_243
timestamp 1649977179
transform 1 0 23460 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_251
timestamp 1649977179
transform 1 0 24196 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_268
timestamp 1649977179
transform 1 0 25760 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_274
timestamp 1649977179
transform 1 0 26312 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_297
timestamp 1649977179
transform 1 0 28428 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_303
timestamp 1649977179
transform 1 0 28980 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_320
timestamp 1649977179
transform 1 0 30544 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1649977179
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_345
timestamp 1649977179
transform 1 0 32844 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_363
timestamp 1649977179
transform 1 0 34500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_375
timestamp 1649977179
transform 1 0 35604 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_384
timestamp 1649977179
transform 1 0 36432 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_395
timestamp 1649977179
transform 1 0 37444 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_401
timestamp 1649977179
transform 1 0 37996 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_124
timestamp 1649977179
transform 1 0 12512 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_136
timestamp 1649977179
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_149
timestamp 1649977179
transform 1 0 14812 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_158
timestamp 1649977179
transform 1 0 15640 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_170
timestamp 1649977179
transform 1 0 16744 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_176
timestamp 1649977179
transform 1 0 17296 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_188
timestamp 1649977179
transform 1 0 18400 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_199
timestamp 1649977179
transform 1 0 19412 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_206
timestamp 1649977179
transform 1 0 20056 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_214
timestamp 1649977179
transform 1 0 20792 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_227
timestamp 1649977179
transform 1 0 21988 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_236
timestamp 1649977179
transform 1 0 22816 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_242
timestamp 1649977179
transform 1 0 23368 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1649977179
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_257
timestamp 1649977179
transform 1 0 24748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_264
timestamp 1649977179
transform 1 0 25392 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_270
timestamp 1649977179
transform 1 0 25944 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_281
timestamp 1649977179
transform 1 0 26956 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_287
timestamp 1649977179
transform 1 0 27508 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_293
timestamp 1649977179
transform 1 0 28060 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_299
timestamp 1649977179
transform 1 0 28612 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_313
timestamp 1649977179
transform 1 0 29900 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_330
timestamp 1649977179
transform 1 0 31464 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_336
timestamp 1649977179
transform 1 0 32016 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_353
timestamp 1649977179
transform 1 0 33580 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_359
timestamp 1649977179
transform 1 0 34132 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_381
timestamp 1649977179
transform 1 0 36156 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_403
timestamp 1649977179
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_77
timestamp 1649977179
transform 1 0 8188 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_82
timestamp 1649977179
transform 1 0 8648 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_90
timestamp 1649977179
transform 1 0 9384 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_94
timestamp 1649977179
transform 1 0 9752 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_106
timestamp 1649977179
transform 1 0 10856 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_139
timestamp 1649977179
transform 1 0 13892 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_145
timestamp 1649977179
transform 1 0 14444 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_154
timestamp 1649977179
transform 1 0 15272 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1649977179
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_173
timestamp 1649977179
transform 1 0 17020 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_176
timestamp 1649977179
transform 1 0 17296 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_180
timestamp 1649977179
transform 1 0 17664 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_183
timestamp 1649977179
transform 1 0 17940 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_187
timestamp 1649977179
transform 1 0 18308 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_190
timestamp 1649977179
transform 1 0 18584 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_203
timestamp 1649977179
transform 1 0 19780 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_210
timestamp 1649977179
transform 1 0 20424 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_218
timestamp 1649977179
transform 1 0 21160 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_234
timestamp 1649977179
transform 1 0 22632 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_247
timestamp 1649977179
transform 1 0 23828 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_267
timestamp 1649977179
transform 1 0 25668 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_274
timestamp 1649977179
transform 1 0 26312 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_284
timestamp 1649977179
transform 1 0 27232 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_290
timestamp 1649977179
transform 1 0 27784 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_310
timestamp 1649977179
transform 1 0 29624 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_316
timestamp 1649977179
transform 1 0 30176 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_322
timestamp 1649977179
transform 1 0 30728 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_328
timestamp 1649977179
transform 1 0 31280 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_339
timestamp 1649977179
transform 1 0 32292 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_343
timestamp 1649977179
transform 1 0 32660 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_348
timestamp 1649977179
transform 1 0 33120 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_356
timestamp 1649977179
transform 1 0 33856 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_364
timestamp 1649977179
transform 1 0 34592 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_370
timestamp 1649977179
transform 1 0 35144 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_376
timestamp 1649977179
transform 1 0 35696 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_384
timestamp 1649977179
transform 1 0 36432 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_397
timestamp 1649977179
transform 1 0 37628 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_402
timestamp 1649977179
transform 1 0 38088 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_406
timestamp 1649977179
transform 1 0 38456 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_18
timestamp 1649977179
transform 1 0 2760 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1649977179
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_35
timestamp 1649977179
transform 1 0 4324 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_38
timestamp 1649977179
transform 1 0 4600 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_44
timestamp 1649977179
transform 1 0 5152 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_50
timestamp 1649977179
transform 1 0 5704 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_58
timestamp 1649977179
transform 1 0 6440 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_63
timestamp 1649977179
transform 1 0 6900 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_69
timestamp 1649977179
transform 1 0 7452 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1649977179
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_89
timestamp 1649977179
transform 1 0 9292 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_92
timestamp 1649977179
transform 1 0 9568 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_62_102
timestamp 1649977179
transform 1 0 10488 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_110
timestamp 1649977179
transform 1 0 11224 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_118
timestamp 1649977179
transform 1 0 11960 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_122
timestamp 1649977179
transform 1 0 12328 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_128
timestamp 1649977179
transform 1 0 12880 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1649977179
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_146
timestamp 1649977179
transform 1 0 14536 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_152
timestamp 1649977179
transform 1 0 15088 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_155
timestamp 1649977179
transform 1 0 15364 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_161
timestamp 1649977179
transform 1 0 15916 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_167
timestamp 1649977179
transform 1 0 16468 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_173
timestamp 1649977179
transform 1 0 17020 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_179
timestamp 1649977179
transform 1 0 17572 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_185
timestamp 1649977179
transform 1 0 18124 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1649977179
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_203
timestamp 1649977179
transform 1 0 19780 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_216
timestamp 1649977179
transform 1 0 20976 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_229
timestamp 1649977179
transform 1 0 22172 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_236
timestamp 1649977179
transform 1 0 22816 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_243
timestamp 1649977179
transform 1 0 23460 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_256
timestamp 1649977179
transform 1 0 24656 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_260
timestamp 1649977179
transform 1 0 25024 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_285
timestamp 1649977179
transform 1 0 27324 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_302
timestamp 1649977179
transform 1 0 28888 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_311
timestamp 1649977179
transform 1 0 29716 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_315
timestamp 1649977179
transform 1 0 30084 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_332
timestamp 1649977179
transform 1 0 31648 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_356
timestamp 1649977179
transform 1 0 33856 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_369
timestamp 1649977179
transform 1 0 35052 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_386
timestamp 1649977179
transform 1 0 36616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_394
timestamp 1649977179
transform 1 0 37352 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_402
timestamp 1649977179
transform 1 0 38088 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_406
timestamp 1649977179
transform 1 0 38456 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_7
timestamp 1649977179
transform 1 0 1748 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_10
timestamp 1649977179
transform 1 0 2024 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_16
timestamp 1649977179
transform 1 0 2576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_22
timestamp 1649977179
transform 1 0 3128 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_30
timestamp 1649977179
transform 1 0 3864 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_42
timestamp 1649977179
transform 1 0 4968 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1649977179
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_61
timestamp 1649977179
transform 1 0 6716 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_67
timestamp 1649977179
transform 1 0 7268 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_70
timestamp 1649977179
transform 1 0 7544 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_78
timestamp 1649977179
transform 1 0 8280 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_90
timestamp 1649977179
transform 1 0 9384 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_100
timestamp 1649977179
transform 1 0 10304 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_108
timestamp 1649977179
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_118
timestamp 1649977179
transform 1 0 11960 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_126
timestamp 1649977179
transform 1 0 12696 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_136
timestamp 1649977179
transform 1 0 13616 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_144
timestamp 1649977179
transform 1 0 14352 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_154
timestamp 1649977179
transform 1 0 15272 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_162
timestamp 1649977179
transform 1 0 16008 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_174
timestamp 1649977179
transform 1 0 17112 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_188
timestamp 1649977179
transform 1 0 18400 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_201
timestamp 1649977179
transform 1 0 19596 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_207
timestamp 1649977179
transform 1 0 20148 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1649977179
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_228
timestamp 1649977179
transform 1 0 22080 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_236
timestamp 1649977179
transform 1 0 22816 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_246
timestamp 1649977179
transform 1 0 23736 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_266
timestamp 1649977179
transform 1 0 25576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1649977179
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_297
timestamp 1649977179
transform 1 0 28428 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_325
timestamp 1649977179
transform 1 0 31004 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_331
timestamp 1649977179
transform 1 0 31556 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_353
timestamp 1649977179
transform 1 0 33580 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_381
timestamp 1649977179
transform 1 0 36156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_387
timestamp 1649977179
transform 1 0 36708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_397
timestamp 1649977179
transform 1 0 37628 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_8
timestamp 1649977179
transform 1 0 1840 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_16
timestamp 1649977179
transform 1 0 2576 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1649977179
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_36
timestamp 1649977179
transform 1 0 4416 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_44
timestamp 1649977179
transform 1 0 5152 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_52
timestamp 1649977179
transform 1 0 5888 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_57
timestamp 1649977179
transform 1 0 6348 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_64
timestamp 1649977179
transform 1 0 6992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_72
timestamp 1649977179
transform 1 0 7728 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_80
timestamp 1649977179
transform 1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_92
timestamp 1649977179
transform 1 0 9568 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_100
timestamp 1649977179
transform 1 0 10304 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_108
timestamp 1649977179
transform 1 0 11040 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_113
timestamp 1649977179
transform 1 0 11500 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_120
timestamp 1649977179
transform 1 0 12144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_128
timestamp 1649977179
transform 1 0 12880 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_136
timestamp 1649977179
transform 1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_148
timestamp 1649977179
transform 1 0 14720 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_156
timestamp 1649977179
transform 1 0 15456 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_164
timestamp 1649977179
transform 1 0 16192 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_169
timestamp 1649977179
transform 1 0 16652 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_173
timestamp 1649977179
transform 1 0 17020 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_178
timestamp 1649977179
transform 1 0 17480 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1649977179
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_204
timestamp 1649977179
transform 1 0 19872 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_211
timestamp 1649977179
transform 1 0 20516 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_218
timestamp 1649977179
transform 1 0 21160 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_228
timestamp 1649977179
transform 1 0 22080 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_235
timestamp 1649977179
transform 1 0 22724 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_242
timestamp 1649977179
transform 1 0 23368 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1649977179
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_256
timestamp 1649977179
transform 1 0 24656 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_263
timestamp 1649977179
transform 1 0 25300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_270
timestamp 1649977179
transform 1 0 25944 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_276
timestamp 1649977179
transform 1 0 26496 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_281
timestamp 1649977179
transform 1 0 26956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_288
timestamp 1649977179
transform 1 0 27600 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_296
timestamp 1649977179
transform 1 0 28336 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1649977179
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_313
timestamp 1649977179
transform 1 0 29900 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_329
timestamp 1649977179
transform 1 0 31372 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1649977179
transform 1 0 31924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_341
timestamp 1649977179
transform 1 0 32476 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_349
timestamp 1649977179
transform 1 0 33212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1649977179
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1649977179
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_367
timestamp 1649977179
transform 1 0 34868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_371
timestamp 1649977179
transform 1 0 35236 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_388
timestamp 1649977179
transform 1 0 36800 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_397
timestamp 1649977179
transform 1 0 37628 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_403
timestamp 1649977179
transform 1 0 38180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_4  _0437_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19320 0 -1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__and2b_1  _0438_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 35880 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0439_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 36340 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0440_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15180 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0441_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15180 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _0442_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16192 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0443_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0444_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15640 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0445_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16376 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0446_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20884 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0447_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17664 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1649977179
transform -1 0 17296 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0449_
timestamp 1649977179
transform 1 0 18492 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0450_
timestamp 1649977179
transform -1 0 21344 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1649977179
transform -1 0 21436 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0452_
timestamp 1649977179
transform -1 0 18492 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0453_
timestamp 1649977179
transform -1 0 18492 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0454_
timestamp 1649977179
transform -1 0 20516 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0455_
timestamp 1649977179
transform -1 0 21620 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0456_
timestamp 1649977179
transform -1 0 21620 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1649977179
transform -1 0 23184 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0458_
timestamp 1649977179
transform -1 0 22632 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1649977179
transform -1 0 22816 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0460_
timestamp 1649977179
transform -1 0 21068 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0461_
timestamp 1649977179
transform -1 0 22080 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0462_
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0463_
timestamp 1649977179
transform 1 0 18768 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0464_
timestamp 1649977179
transform -1 0 18400 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0465_
timestamp 1649977179
transform -1 0 21344 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0466_
timestamp 1649977179
transform -1 0 22080 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0467_
timestamp 1649977179
transform -1 0 22172 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0468_
timestamp 1649977179
transform -1 0 23460 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0469_
timestamp 1649977179
transform -1 0 23828 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1649977179
transform -1 0 24656 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0471_
timestamp 1649977179
transform -1 0 23736 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0472_
timestamp 1649977179
transform -1 0 24656 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0473_
timestamp 1649977179
transform -1 0 22632 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0474_
timestamp 1649977179
transform -1 0 22816 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0475_
timestamp 1649977179
transform 1 0 23000 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0476_
timestamp 1649977179
transform -1 0 22816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0477_
timestamp 1649977179
transform 1 0 22908 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0478_
timestamp 1649977179
transform -1 0 23460 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0479_
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0480_
timestamp 1649977179
transform -1 0 22264 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0481_
timestamp 1649977179
transform -1 0 19780 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0482_
timestamp 1649977179
transform -1 0 20056 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0483_
timestamp 1649977179
transform 1 0 20148 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0484_
timestamp 1649977179
transform -1 0 20516 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13524 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0486_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13892 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0487_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18768 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0488_
timestamp 1649977179
transform -1 0 19964 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1649977179
transform 1 0 11592 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0490_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0491_
timestamp 1649977179
transform 1 0 19044 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0492_
timestamp 1649977179
transform -1 0 20332 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0493_
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0494_
timestamp 1649977179
transform 1 0 18032 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0495_
timestamp 1649977179
transform -1 0 20700 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0496_
timestamp 1649977179
transform 1 0 20516 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0497_
timestamp 1649977179
transform -1 0 22264 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _0498_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16008 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0499_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14444 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _0500_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13892 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0501_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13524 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0502_
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0503_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18400 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0504_
timestamp 1649977179
transform -1 0 13156 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0505_
timestamp 1649977179
transform -1 0 13248 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0506_
timestamp 1649977179
transform -1 0 9568 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0507_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10396 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_2  _0508_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0509_
timestamp 1649977179
transform 1 0 9200 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0510_
timestamp 1649977179
transform -1 0 10672 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0511_
timestamp 1649977179
transform 1 0 10028 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0512_
timestamp 1649977179
transform -1 0 14996 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0513_
timestamp 1649977179
transform 1 0 15364 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0514_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15272 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1649977179
transform -1 0 12880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0516_
timestamp 1649977179
transform 1 0 11960 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _0517_
timestamp 1649977179
transform -1 0 13892 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0518_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14996 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0519_
timestamp 1649977179
transform -1 0 16928 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1649977179
transform -1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0521_
timestamp 1649977179
transform 1 0 13616 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0522_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14168 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0523_
timestamp 1649977179
transform -1 0 16744 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0524_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15456 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0525_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18492 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0526_
timestamp 1649977179
transform -1 0 18216 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_4  _0527_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17204 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_4  _0528_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13064 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0529_
timestamp 1649977179
transform 1 0 12696 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0530_
timestamp 1649977179
transform -1 0 13156 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0531_
timestamp 1649977179
transform 1 0 13524 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0532_
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0533_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0534_
timestamp 1649977179
transform -1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0535_
timestamp 1649977179
transform 1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0536_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0537_
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0538_
timestamp 1649977179
transform -1 0 13156 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0539_
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0540_
timestamp 1649977179
transform 1 0 10028 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0541_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12880 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0542_
timestamp 1649977179
transform -1 0 16192 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0543_
timestamp 1649977179
transform -1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0544_
timestamp 1649977179
transform -1 0 15180 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0545_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0546_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14168 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0547_
timestamp 1649977179
transform -1 0 15916 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0548_
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0549_
timestamp 1649977179
transform -1 0 21528 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0550_
timestamp 1649977179
transform 1 0 20516 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0551_
timestamp 1649977179
transform 1 0 16376 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0552_
timestamp 1649977179
transform -1 0 17480 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0553_
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0554_
timestamp 1649977179
transform -1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0555_
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0556_
timestamp 1649977179
transform -1 0 30360 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0557_
timestamp 1649977179
transform -1 0 17112 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0558_
timestamp 1649977179
transform 1 0 32384 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0559_
timestamp 1649977179
transform -1 0 33488 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0560_
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1649977179
transform -1 0 37996 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0562_
timestamp 1649977179
transform -1 0 22172 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0563_
timestamp 1649977179
transform -1 0 21436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _0564_
timestamp 1649977179
transform 1 0 19780 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0565_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0566_
timestamp 1649977179
transform -1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0567_
timestamp 1649977179
transform -1 0 20056 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0568_
timestamp 1649977179
transform -1 0 20976 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0569_
timestamp 1649977179
transform -1 0 36984 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0570_
timestamp 1649977179
transform -1 0 37536 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0571_
timestamp 1649977179
transform 1 0 36524 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1649977179
transform 1 0 36248 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0573_
timestamp 1649977179
transform 1 0 16744 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0574_
timestamp 1649977179
transform -1 0 34316 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0575_
timestamp 1649977179
transform -1 0 34960 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0576_
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0577_
timestamp 1649977179
transform -1 0 18400 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0578_
timestamp 1649977179
transform -1 0 17480 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1649977179
transform -1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0580_
timestamp 1649977179
transform -1 0 18400 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1649977179
transform -1 0 24840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0582_
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0583_
timestamp 1649977179
transform 1 0 29900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0584_
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0585_
timestamp 1649977179
transform -1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0586_
timestamp 1649977179
transform -1 0 31280 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0587_
timestamp 1649977179
transform -1 0 32384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0588_
timestamp 1649977179
transform -1 0 32936 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0589_
timestamp 1649977179
transform -1 0 34224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0590_
timestamp 1649977179
transform -1 0 34224 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0591_
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0592_
timestamp 1649977179
transform -1 0 31924 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0593_
timestamp 1649977179
transform 1 0 37444 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0594_
timestamp 1649977179
transform 1 0 19596 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0595_
timestamp 1649977179
transform -1 0 33304 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0596_
timestamp 1649977179
transform -1 0 36248 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0597_
timestamp 1649977179
transform -1 0 34224 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0598_
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0599_
timestamp 1649977179
transform -1 0 35512 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0600_
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0601_
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0602_
timestamp 1649977179
transform -1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0603_
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0604_
timestamp 1649977179
transform -1 0 34960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0605_
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0606_
timestamp 1649977179
transform -1 0 34224 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0607_
timestamp 1649977179
transform -1 0 34868 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1649977179
transform -1 0 36340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0609_
timestamp 1649977179
transform -1 0 20056 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0610_
timestamp 1649977179
transform -1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0611_
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0612_
timestamp 1649977179
transform -1 0 19136 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0613_
timestamp 1649977179
transform -1 0 20056 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0614_
timestamp 1649977179
transform -1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0615_
timestamp 1649977179
transform -1 0 11040 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0616_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0617_
timestamp 1649977179
transform -1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0618_
timestamp 1649977179
transform -1 0 10764 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0619_
timestamp 1649977179
transform -1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0620_
timestamp 1649977179
transform -1 0 11040 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1649977179
transform -1 0 11776 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1649977179
transform -1 0 10028 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0623_
timestamp 1649977179
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0624_
timestamp 1649977179
transform -1 0 9660 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0625_
timestamp 1649977179
transform -1 0 9384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0626_
timestamp 1649977179
transform -1 0 12512 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0627_
timestamp 1649977179
transform -1 0 13432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0628_
timestamp 1649977179
transform -1 0 12328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0629_
timestamp 1649977179
transform -1 0 12144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0630_
timestamp 1649977179
transform -1 0 11040 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0631_
timestamp 1649977179
transform -1 0 11132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0632_
timestamp 1649977179
transform -1 0 10672 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1649977179
transform -1 0 10672 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0634_
timestamp 1649977179
transform -1 0 12420 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0635_
timestamp 1649977179
transform -1 0 13248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0636_
timestamp 1649977179
transform 1 0 14628 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0637_
timestamp 1649977179
transform -1 0 15916 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0638_
timestamp 1649977179
transform -1 0 15824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0639_
timestamp 1649977179
transform 1 0 14168 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0640_
timestamp 1649977179
transform -1 0 14628 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0641_
timestamp 1649977179
transform 1 0 13892 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1649977179
transform -1 0 13616 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0643_
timestamp 1649977179
transform 1 0 13892 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 1649977179
transform -1 0 14352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0645_
timestamp 1649977179
transform -1 0 16008 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0646_
timestamp 1649977179
transform -1 0 16192 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0647_
timestamp 1649977179
transform -1 0 17480 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1649977179
transform -1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0649_
timestamp 1649977179
transform -1 0 17388 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0650_
timestamp 1649977179
transform -1 0 19688 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0651_
timestamp 1649977179
transform -1 0 17572 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0652_
timestamp 1649977179
transform -1 0 18400 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0653_
timestamp 1649977179
transform 1 0 18124 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1649977179
transform -1 0 17756 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0655_
timestamp 1649977179
transform -1 0 18400 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0656_
timestamp 1649977179
transform -1 0 18308 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0657_
timestamp 1649977179
transform -1 0 20148 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0658_
timestamp 1649977179
transform -1 0 20700 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0659_
timestamp 1649977179
transform -1 0 18768 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1649977179
transform -1 0 18768 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0661_
timestamp 1649977179
transform -1 0 29072 0 1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_4  _0662_
timestamp 1649977179
transform -1 0 20700 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0663_
timestamp 1649977179
transform 1 0 16468 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0664_
timestamp 1649977179
transform 1 0 15272 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0665_
timestamp 1649977179
transform -1 0 16928 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0666_
timestamp 1649977179
transform 1 0 17204 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0667_
timestamp 1649977179
transform 1 0 15732 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0668_
timestamp 1649977179
transform -1 0 17756 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0669_
timestamp 1649977179
transform 1 0 17756 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0670_
timestamp 1649977179
transform 1 0 16560 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0671_
timestamp 1649977179
transform -1 0 18124 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0672_
timestamp 1649977179
transform 1 0 16560 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0673_
timestamp 1649977179
transform 1 0 15916 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0674_
timestamp 1649977179
transform -1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0675_
timestamp 1649977179
transform 1 0 17940 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0676_
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0677_
timestamp 1649977179
transform -1 0 17480 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0678_
timestamp 1649977179
transform 1 0 20516 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0679_
timestamp 1649977179
transform 1 0 17480 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0680_
timestamp 1649977179
transform -1 0 18492 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0681_
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0682_
timestamp 1649977179
transform 1 0 17848 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0683_
timestamp 1649977179
transform -1 0 19504 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0684_
timestamp 1649977179
transform -1 0 19596 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0685_
timestamp 1649977179
transform -1 0 19688 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0686_
timestamp 1649977179
transform -1 0 18768 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0687_
timestamp 1649977179
transform 1 0 19412 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0688_
timestamp 1649977179
transform 1 0 18768 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0689_
timestamp 1649977179
transform -1 0 19504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0690_
timestamp 1649977179
transform 1 0 19780 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0691_
timestamp 1649977179
transform 1 0 19688 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0692_
timestamp 1649977179
transform -1 0 20792 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0693_
timestamp 1649977179
transform 1 0 19964 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0694_
timestamp 1649977179
transform 1 0 19596 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0695_
timestamp 1649977179
transform -1 0 20332 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0696_
timestamp 1649977179
transform 1 0 21712 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0697_
timestamp 1649977179
transform -1 0 20884 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0698_
timestamp 1649977179
transform -1 0 19780 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0699_
timestamp 1649977179
transform 1 0 20056 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0700_
timestamp 1649977179
transform -1 0 20424 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0701_
timestamp 1649977179
transform -1 0 20148 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0702_
timestamp 1649977179
transform -1 0 21804 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0703_
timestamp 1649977179
transform -1 0 22264 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0704_
timestamp 1649977179
transform -1 0 21988 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0705_
timestamp 1649977179
transform 1 0 22724 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0706_
timestamp 1649977179
transform 1 0 22356 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0707_
timestamp 1649977179
transform -1 0 23460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0708_
timestamp 1649977179
transform 1 0 24472 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0709_
timestamp 1649977179
transform 1 0 23460 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0710_
timestamp 1649977179
transform -1 0 24656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0711_
timestamp 1649977179
transform -1 0 25392 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0712_
timestamp 1649977179
transform 1 0 26036 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0713_
timestamp 1649977179
transform -1 0 28796 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0714_
timestamp 1649977179
transform -1 0 25944 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0715_
timestamp 1649977179
transform 1 0 26220 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0716_
timestamp 1649977179
transform -1 0 30544 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0717_
timestamp 1649977179
transform 1 0 23368 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0718_
timestamp 1649977179
transform -1 0 28152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0719_
timestamp 1649977179
transform 1 0 31740 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0720_
timestamp 1649977179
transform -1 0 33304 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0721_
timestamp 1649977179
transform -1 0 29992 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0722_
timestamp 1649977179
transform -1 0 29808 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0723_
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0724_
timestamp 1649977179
transform 1 0 17480 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0725_
timestamp 1649977179
transform -1 0 22448 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0726_
timestamp 1649977179
transform -1 0 20884 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0727_
timestamp 1649977179
transform 1 0 20792 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0728_
timestamp 1649977179
transform 1 0 25576 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0729_
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0730_
timestamp 1649977179
transform -1 0 24840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0731_
timestamp 1649977179
transform 1 0 22172 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0732_
timestamp 1649977179
transform 1 0 22172 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0733_
timestamp 1649977179
transform -1 0 23368 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0734_
timestamp 1649977179
transform 1 0 22080 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0735_
timestamp 1649977179
transform 1 0 21896 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0736_
timestamp 1649977179
transform -1 0 22724 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0737_
timestamp 1649977179
transform 1 0 35512 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0738_
timestamp 1649977179
transform 1 0 29624 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0739_
timestamp 1649977179
transform -1 0 31280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0740_
timestamp 1649977179
transform 1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0741_
timestamp 1649977179
transform 1 0 36064 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0742_
timestamp 1649977179
transform 1 0 36064 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0743_
timestamp 1649977179
transform 1 0 36800 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 1649977179
transform -1 0 38180 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0745_
timestamp 1649977179
transform 1 0 37720 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0746_
timestamp 1649977179
transform 1 0 37812 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0747_
timestamp 1649977179
transform -1 0 22632 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0748_
timestamp 1649977179
transform 1 0 23000 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0749_
timestamp 1649977179
transform -1 0 25484 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0750_
timestamp 1649977179
transform 1 0 26128 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0751_
timestamp 1649977179
transform 1 0 25392 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0752_
timestamp 1649977179
transform -1 0 27324 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0753_
timestamp 1649977179
transform 1 0 28336 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0754_
timestamp 1649977179
transform -1 0 28520 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0755_
timestamp 1649977179
transform -1 0 27968 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 1649977179
transform -1 0 28704 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0757_
timestamp 1649977179
transform -1 0 28888 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0758_
timestamp 1649977179
transform -1 0 28612 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0759_
timestamp 1649977179
transform 1 0 21712 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 1649977179
transform 1 0 27968 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0761_
timestamp 1649977179
transform 1 0 27600 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0762_
timestamp 1649977179
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0763_
timestamp 1649977179
transform 1 0 29532 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0764_
timestamp 1649977179
transform 1 0 29624 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0765_
timestamp 1649977179
transform -1 0 30636 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0766_
timestamp 1649977179
transform 1 0 30912 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0767_
timestamp 1649977179
transform 1 0 30728 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0768_
timestamp 1649977179
transform -1 0 31832 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0769_
timestamp 1649977179
transform 1 0 29716 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0770_
timestamp 1649977179
transform 1 0 29808 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0771_
timestamp 1649977179
transform -1 0 32384 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0772_
timestamp 1649977179
transform 1 0 18952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0773_
timestamp 1649977179
transform 1 0 30820 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0774_
timestamp 1649977179
transform 1 0 30820 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0775_
timestamp 1649977179
transform -1 0 31464 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0776_
timestamp 1649977179
transform 1 0 33396 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0777_
timestamp 1649977179
transform 1 0 32936 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0778_
timestamp 1649977179
transform -1 0 36248 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0779_
timestamp 1649977179
transform 1 0 35696 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0780_
timestamp 1649977179
transform -1 0 35788 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0781_
timestamp 1649977179
transform -1 0 35604 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0783_
timestamp 1649977179
transform -1 0 34316 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0784_
timestamp 1649977179
transform -1 0 33948 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1649977179
transform 1 0 35880 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0786_
timestamp 1649977179
transform -1 0 35972 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0787_
timestamp 1649977179
transform 1 0 35512 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1649977179
transform 1 0 35236 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0789_
timestamp 1649977179
transform -1 0 35144 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0790_
timestamp 1649977179
transform -1 0 34960 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0791_
timestamp 1649977179
transform -1 0 19964 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 1649977179
transform 1 0 32752 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0793_
timestamp 1649977179
transform 1 0 32476 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0794_
timestamp 1649977179
transform -1 0 35420 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 1649977179
transform -1 0 34868 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0796_
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0797_
timestamp 1649977179
transform -1 0 36616 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0798_
timestamp 1649977179
transform -1 0 20056 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0799_
timestamp 1649977179
transform 1 0 19596 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0800_
timestamp 1649977179
transform -1 0 21252 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1649977179
transform -1 0 18676 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0802_
timestamp 1649977179
transform 1 0 18308 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0803_
timestamp 1649977179
transform -1 0 18952 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0804_
timestamp 1649977179
transform -1 0 14536 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1649977179
transform -1 0 14904 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0806_
timestamp 1649977179
transform 1 0 14352 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0807_
timestamp 1649977179
transform -1 0 14996 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1649977179
transform 1 0 10212 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0809_
timestamp 1649977179
transform 1 0 10396 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0810_
timestamp 1649977179
transform -1 0 11960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0811_
timestamp 1649977179
transform 1 0 9016 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0812_
timestamp 1649977179
transform 1 0 8832 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0813_
timestamp 1649977179
transform -1 0 10028 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0815_
timestamp 1649977179
transform 1 0 8372 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0816_
timestamp 1649977179
transform -1 0 9384 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0817_
timestamp 1649977179
transform 1 0 9108 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0818_
timestamp 1649977179
transform 1 0 9200 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0819_
timestamp 1649977179
transform -1 0 10304 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0820_
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0821_
timestamp 1649977179
transform 1 0 10856 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0822_
timestamp 1649977179
transform -1 0 11868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0823_
timestamp 1649977179
transform -1 0 17572 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0824_
timestamp 1649977179
transform 1 0 12328 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0825_
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0826_
timestamp 1649977179
transform -1 0 12880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0827_
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0828_
timestamp 1649977179
transform 1 0 11776 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0829_
timestamp 1649977179
transform -1 0 12512 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0830_
timestamp 1649977179
transform 1 0 11960 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0831_
timestamp 1649977179
transform 1 0 11868 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0832_
timestamp 1649977179
transform -1 0 12420 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0833_
timestamp 1649977179
transform 1 0 11592 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0834_
timestamp 1649977179
transform 1 0 10856 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0835_
timestamp 1649977179
transform -1 0 11868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0836_
timestamp 1649977179
transform 1 0 14904 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0837_
timestamp 1649977179
transform 1 0 13248 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0838_
timestamp 1649977179
transform -1 0 13156 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0839_
timestamp 1649977179
transform -1 0 13248 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0840_
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0841_
timestamp 1649977179
transform 1 0 15180 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0842_
timestamp 1649977179
transform -1 0 16928 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0843_
timestamp 1649977179
transform 1 0 15364 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0844_
timestamp 1649977179
transform 1 0 15088 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0845_
timestamp 1649977179
transform -1 0 16928 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0846_
timestamp 1649977179
transform 1 0 14444 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0847_
timestamp 1649977179
transform -1 0 14536 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0848_
timestamp 1649977179
transform -1 0 14352 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0849_
timestamp 1649977179
transform -1 0 15916 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0850_
timestamp 1649977179
transform 1 0 15272 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0851_
timestamp 1649977179
transform -1 0 16928 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0852_
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0853_
timestamp 1649977179
transform 1 0 16744 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0854_
timestamp 1649977179
transform -1 0 18124 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0855_
timestamp 1649977179
transform 1 0 17204 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0856_
timestamp 1649977179
transform 1 0 17020 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0857_
timestamp 1649977179
transform -1 0 17756 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 1649977179
transform -1 0 17480 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0859_
timestamp 1649977179
transform 1 0 17388 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0860_
timestamp 1649977179
transform -1 0 18768 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0861_
timestamp 1649977179
transform -1 0 18768 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0862_
timestamp 1649977179
transform 1 0 18768 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0863_
timestamp 1649977179
transform -1 0 19780 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0864_
timestamp 1649977179
transform 1 0 19596 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0865_
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0866_
timestamp 1649977179
transform -1 0 19964 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0867_
timestamp 1649977179
transform 1 0 21160 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0868_
timestamp 1649977179
transform 1 0 20424 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0869_
timestamp 1649977179
transform -1 0 21896 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0870_
timestamp 1649977179
transform -1 0 20884 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0871_
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0872_
timestamp 1649977179
transform -1 0 22540 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0873_
timestamp 1649977179
transform -1 0 21160 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0874_
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0875_
timestamp 1649977179
transform -1 0 22908 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0876_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24472 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0877_
timestamp 1649977179
transform -1 0 26496 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0878_
timestamp 1649977179
transform -1 0 29072 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0879_
timestamp 1649977179
transform -1 0 31924 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0880_
timestamp 1649977179
transform 1 0 26864 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0881_
timestamp 1649977179
transform -1 0 25760 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0882_
timestamp 1649977179
transform -1 0 25852 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0883_
timestamp 1649977179
transform 1 0 29992 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0884_
timestamp 1649977179
transform -1 0 25576 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0885_
timestamp 1649977179
transform -1 0 30268 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0886_
timestamp 1649977179
transform -1 0 28428 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0887_
timestamp 1649977179
transform 1 0 30176 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0888_
timestamp 1649977179
transform -1 0 33580 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0889_
timestamp 1649977179
transform -1 0 28888 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0890_
timestamp 1649977179
transform -1 0 29624 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0891_
timestamp 1649977179
transform -1 0 33856 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0892_
timestamp 1649977179
transform -1 0 34500 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0893_
timestamp 1649977179
transform -1 0 36156 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0894_
timestamp 1649977179
transform -1 0 35420 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0895_
timestamp 1649977179
transform -1 0 33764 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0896_
timestamp 1649977179
transform -1 0 30728 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0897_
timestamp 1649977179
transform -1 0 25852 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0898_
timestamp 1649977179
transform -1 0 29256 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0899_
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0900_
timestamp 1649977179
transform -1 0 28152 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0901_
timestamp 1649977179
transform -1 0 30544 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0902_
timestamp 1649977179
transform -1 0 26588 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0903_
timestamp 1649977179
transform -1 0 25668 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0904_
timestamp 1649977179
transform -1 0 23552 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0905_
timestamp 1649977179
transform -1 0 28428 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0906_
timestamp 1649977179
transform -1 0 23736 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0907_
timestamp 1649977179
transform -1 0 28520 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0908_
timestamp 1649977179
transform -1 0 26680 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0909_
timestamp 1649977179
transform -1 0 31004 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0910_
timestamp 1649977179
transform -1 0 30268 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0911_
timestamp 1649977179
transform -1 0 36156 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0912_
timestamp 1649977179
transform -1 0 33580 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0913_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 38180 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0914_
timestamp 1649977179
transform -1 0 30544 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0915_
timestamp 1649977179
transform -1 0 28428 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0916_
timestamp 1649977179
transform -1 0 25116 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0917_
timestamp 1649977179
transform -1 0 23276 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0918_
timestamp 1649977179
transform -1 0 38180 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0919_
timestamp 1649977179
transform 1 0 36064 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0920_
timestamp 1649977179
transform -1 0 35420 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0921_
timestamp 1649977179
transform -1 0 28428 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0922_
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0923_
timestamp 1649977179
transform 1 0 27048 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0924_
timestamp 1649977179
transform 1 0 29532 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0925_
timestamp 1649977179
transform 1 0 32384 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0926_
timestamp 1649977179
transform -1 0 33120 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0927_
timestamp 1649977179
transform 1 0 36156 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0928_
timestamp 1649977179
transform 1 0 32568 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0929_
timestamp 1649977179
transform -1 0 36800 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0930_
timestamp 1649977179
transform 1 0 35972 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0931_
timestamp 1649977179
transform -1 0 36524 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0932_
timestamp 1649977179
transform -1 0 36800 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0933_
timestamp 1649977179
transform 1 0 36708 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0934_
timestamp 1649977179
transform 1 0 34868 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0935_
timestamp 1649977179
transform -1 0 37076 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0936_
timestamp 1649977179
transform 1 0 36708 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0937_
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0938_
timestamp 1649977179
transform -1 0 29900 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0939_
timestamp 1649977179
transform 1 0 21344 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0940_
timestamp 1649977179
transform -1 0 26680 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0941_
timestamp 1649977179
transform -1 0 25484 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0942_
timestamp 1649977179
transform -1 0 27232 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0943_
timestamp 1649977179
transform -1 0 23184 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0944_
timestamp 1649977179
transform 1 0 24104 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0945_
timestamp 1649977179
transform -1 0 23000 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0946_
timestamp 1649977179
transform -1 0 23092 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0947_
timestamp 1649977179
transform -1 0 23276 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0948_
timestamp 1649977179
transform -1 0 23092 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0949_
timestamp 1649977179
transform 1 0 24472 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0950_
timestamp 1649977179
transform -1 0 23276 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0951_
timestamp 1649977179
transform -1 0 25944 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0952_
timestamp 1649977179
transform -1 0 23092 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0953_
timestamp 1649977179
transform -1 0 23276 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0954_
timestamp 1649977179
transform -1 0 23184 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0955_
timestamp 1649977179
transform 1 0 25024 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0956_
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0957_
timestamp 1649977179
transform -1 0 23092 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0958_
timestamp 1649977179
transform -1 0 25576 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0959_
timestamp 1649977179
transform -1 0 28520 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0960_
timestamp 1649977179
transform -1 0 23276 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0961_
timestamp 1649977179
transform -1 0 27692 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0962_
timestamp 1649977179
transform -1 0 27232 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0963_
timestamp 1649977179
transform -1 0 29072 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0964_
timestamp 1649977179
transform -1 0 31832 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0965_
timestamp 1649977179
transform -1 0 31004 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0966_
timestamp 1649977179
transform -1 0 28336 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 1649977179
transform -1 0 28980 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 1649977179
transform -1 0 27784 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0969_
timestamp 1649977179
transform -1 0 28428 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0970_
timestamp 1649977179
transform -1 0 28888 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0971_
timestamp 1649977179
transform -1 0 32016 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1649977179
transform -1 0 36432 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1649977179
transform 1 0 28520 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0974_
timestamp 1649977179
transform -1 0 30820 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1649977179
transform -1 0 33672 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0976_
timestamp 1649977179
transform -1 0 34500 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0977_
timestamp 1649977179
transform 1 0 32200 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1649977179
transform -1 0 32660 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1649977179
transform -1 0 31188 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1649977179
transform -1 0 35512 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1649977179
transform -1 0 34960 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1649977179
transform -1 0 30084 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1649977179
transform 1 0 22172 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1649977179
transform 1 0 28888 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0985_
timestamp 1649977179
transform -1 0 27784 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0986_
timestamp 1649977179
transform 1 0 29716 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1649977179
transform 1 0 35328 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1649977179
transform 1 0 35144 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1649977179
transform 1 0 36708 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1649977179
transform -1 0 32108 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1649977179
transform -1 0 34224 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1649977179
transform -1 0 37076 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1649977179
transform -1 0 34316 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1649977179
transform -1 0 33580 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1649977179
transform -1 0 32384 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1649977179
transform -1 0 33580 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1649977179
transform 1 0 36708 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1649977179
transform 1 0 36708 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1649977179
transform 1 0 36708 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1649977179
transform 1 0 35328 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1649977179
transform 1 0 33948 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1649977179
transform 1 0 34868 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1649977179
transform 1 0 35052 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1649977179
transform 1 0 36708 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1649977179
transform 1 0 36708 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1649977179
transform -1 0 29164 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1649977179
transform -1 0 27692 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1649977179
transform -1 0 25852 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1649977179
transform -1 0 28428 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1649977179
transform -1 0 25852 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1649977179
transform -1 0 25852 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1649977179
transform -1 0 25576 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1649977179
transform -1 0 25852 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1649977179
transform -1 0 25852 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1649977179
transform -1 0 26128 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1649977179
transform -1 0 28520 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1649977179
transform -1 0 25484 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1649977179
transform -1 0 25852 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1649977179
transform -1 0 25760 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1649977179
transform -1 0 28428 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1649977179
transform 1 0 29624 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1649977179
transform 1 0 34684 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1649977179
transform -1 0 32752 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1649977179
transform -1 0 32384 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1649977179
transform -1 0 29440 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1649977179
transform -1 0 33580 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1649977179
transform -1 0 32844 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1649977179
transform 1 0 34960 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_m opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 32016 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_s
timestamp 1649977179
transform -1 0 34316 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk_m
timestamp 1649977179
transform -1 0 25208 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk_s
timestamp 1649977179
transform -1 0 27876 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk_m
timestamp 1649977179
transform -1 0 27876 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk_s
timestamp 1649977179
transform -1 0 30452 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk_m
timestamp 1649977179
transform -1 0 25208 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk_s
timestamp 1649977179
transform -1 0 27876 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk_m
timestamp 1649977179
transform 1 0 26036 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk_s
timestamp 1649977179
transform 1 0 28612 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk_m
timestamp 1649977179
transform -1 0 33028 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk_s
timestamp 1649977179
transform 1 0 31188 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk_m
timestamp 1649977179
transform 1 0 33764 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk_s
timestamp 1649977179
transform 1 0 36340 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk_m
timestamp 1649977179
transform 1 0 31188 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk_s
timestamp 1649977179
transform -1 0 33028 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk_m
timestamp 1649977179
transform 1 0 33764 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk_s
timestamp 1649977179
transform 1 0 33764 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1649977179
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2392 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 11776 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 12972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 4600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform -1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 5888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 7820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform -1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform 1 0 28244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform -1 0 33212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform -1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform -1 0 34224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform 1 0 37444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform 1 0 37904 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform 1 0 35972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 30452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 30912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform 1 0 33948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform -1 0 31648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform 1 0 32292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform 1 0 36800 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 37904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1649977179
transform 1 0 37904 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input48
timestamp 1649977179
transform -1 0 38180 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform 1 0 1472 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform 1 0 3496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1649977179
transform 1 0 17848 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1649977179
transform -1 0 17756 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform 1 0 25944 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform 1 0 24472 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform 1 0 25116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform 1 0 26036 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform 1 0 26680 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1649977179
transform -1 0 18768 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform -1 0 20424 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform -1 0 19872 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform 1 0 20884 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1649977179
transform 1 0 21804 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1649977179
transform 1 0 22448 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1649977179
transform 1 0 23092 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1649977179
transform 1 0 25024 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1649977179
transform 1 0 25668 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform 1 0 16928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 24748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 26220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 25484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 28796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 20792 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 20976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform -1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 24012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform -1 0 23552 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 2576 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform -1 0 4416 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform -1 0 9568 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform -1 0 10304 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform 1 0 10672 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 12144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 12696 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 12512 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 14352 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 14720 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 4968 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 15456 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 16008 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform 1 0 15824 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 17112 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform -1 0 5152 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform -1 0 5888 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform -1 0 6716 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform -1 0 6992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform -1 0 7728 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform -1 0 8280 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform -1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform -1 0 9384 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform -1 0 17480 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform -1 0 27600 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform -1 0 33120 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform -1 0 33856 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform -1 0 34592 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform -1 0 36156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1649977179
transform -1 0 37628 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform -1 0 37628 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform -1 0 28336 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform -1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform -1 0 29900 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform -1 0 30636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform -1 0 31372 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform -1 0 31004 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform -1 0 32476 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform -1 0 33212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform -1 0 33948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform -1 0 36432 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform 1 0 36984 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform 1 0 37720 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform -1 0 38088 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  wb_cross_clk_132 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15916 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 clk_m
port 0 nsew signal input
flabel metal2 s 38198 39200 38254 40000 0 FreeSans 224 90 0 0 clk_s
port 1 nsew signal input
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 m_rst
port 2 nsew signal input
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 m_wb_4_burst
port 3 nsew signal input
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 m_wb_8_burst
port 4 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 m_wb_ack
port 5 nsew signal tristate
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 m_wb_adr[0]
port 6 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 m_wb_adr[10]
port 7 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 m_wb_adr[11]
port 8 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 m_wb_adr[12]
port 9 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 m_wb_adr[13]
port 10 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 m_wb_adr[14]
port 11 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 m_wb_adr[15]
port 12 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 m_wb_adr[16]
port 13 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 m_wb_adr[17]
port 14 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 m_wb_adr[18]
port 15 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 m_wb_adr[19]
port 16 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 m_wb_adr[1]
port 17 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 m_wb_adr[20]
port 18 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 m_wb_adr[21]
port 19 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 m_wb_adr[22]
port 20 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 m_wb_adr[23]
port 21 nsew signal input
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 m_wb_adr[2]
port 22 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 m_wb_adr[3]
port 23 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 m_wb_adr[4]
port 24 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 m_wb_adr[5]
port 25 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 m_wb_adr[6]
port 26 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 m_wb_adr[7]
port 27 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 m_wb_adr[8]
port 28 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 m_wb_adr[9]
port 29 nsew signal input
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 m_wb_cyc
port 30 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 m_wb_err
port 31 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 m_wb_i_dat[0]
port 32 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 m_wb_i_dat[10]
port 33 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 m_wb_i_dat[11]
port 34 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 m_wb_i_dat[12]
port 35 nsew signal tristate
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 m_wb_i_dat[13]
port 36 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 m_wb_i_dat[14]
port 37 nsew signal tristate
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 m_wb_i_dat[15]
port 38 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 m_wb_i_dat[1]
port 39 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 m_wb_i_dat[2]
port 40 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 m_wb_i_dat[3]
port 41 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 m_wb_i_dat[4]
port 42 nsew signal tristate
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 m_wb_i_dat[5]
port 43 nsew signal tristate
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 m_wb_i_dat[6]
port 44 nsew signal tristate
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 m_wb_i_dat[7]
port 45 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 m_wb_i_dat[8]
port 46 nsew signal tristate
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 m_wb_i_dat[9]
port 47 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 m_wb_o_dat[0]
port 48 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 m_wb_o_dat[10]
port 49 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 m_wb_o_dat[11]
port 50 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 m_wb_o_dat[12]
port 51 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 m_wb_o_dat[13]
port 52 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 m_wb_o_dat[14]
port 53 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 m_wb_o_dat[15]
port 54 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 m_wb_o_dat[1]
port 55 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 m_wb_o_dat[2]
port 56 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 m_wb_o_dat[3]
port 57 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 m_wb_o_dat[4]
port 58 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 m_wb_o_dat[5]
port 59 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 m_wb_o_dat[6]
port 60 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 m_wb_o_dat[7]
port 61 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 m_wb_o_dat[8]
port 62 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 m_wb_o_dat[9]
port 63 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 m_wb_sel[0]
port 64 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 m_wb_sel[1]
port 65 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 m_wb_stb
port 66 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 m_wb_we
port 67 nsew signal input
flabel metal2 s 1766 39200 1822 40000 0 FreeSans 224 90 0 0 s_rst
port 68 nsew signal input
flabel metal2 s 2318 39200 2374 40000 0 FreeSans 224 90 0 0 s_wb_4_burst
port 69 nsew signal tristate
flabel metal2 s 2870 39200 2926 40000 0 FreeSans 224 90 0 0 s_wb_8_burst
port 70 nsew signal tristate
flabel metal2 s 3422 39200 3478 40000 0 FreeSans 224 90 0 0 s_wb_ack
port 71 nsew signal input
flabel metal2 s 3974 39200 4030 40000 0 FreeSans 224 90 0 0 s_wb_adr[0]
port 72 nsew signal tristate
flabel metal2 s 9494 39200 9550 40000 0 FreeSans 224 90 0 0 s_wb_adr[10]
port 73 nsew signal tristate
flabel metal2 s 10046 39200 10102 40000 0 FreeSans 224 90 0 0 s_wb_adr[11]
port 74 nsew signal tristate
flabel metal2 s 10598 39200 10654 40000 0 FreeSans 224 90 0 0 s_wb_adr[12]
port 75 nsew signal tristate
flabel metal2 s 11150 39200 11206 40000 0 FreeSans 224 90 0 0 s_wb_adr[13]
port 76 nsew signal tristate
flabel metal2 s 11702 39200 11758 40000 0 FreeSans 224 90 0 0 s_wb_adr[14]
port 77 nsew signal tristate
flabel metal2 s 12254 39200 12310 40000 0 FreeSans 224 90 0 0 s_wb_adr[15]
port 78 nsew signal tristate
flabel metal2 s 12806 39200 12862 40000 0 FreeSans 224 90 0 0 s_wb_adr[16]
port 79 nsew signal tristate
flabel metal2 s 13358 39200 13414 40000 0 FreeSans 224 90 0 0 s_wb_adr[17]
port 80 nsew signal tristate
flabel metal2 s 13910 39200 13966 40000 0 FreeSans 224 90 0 0 s_wb_adr[18]
port 81 nsew signal tristate
flabel metal2 s 14462 39200 14518 40000 0 FreeSans 224 90 0 0 s_wb_adr[19]
port 82 nsew signal tristate
flabel metal2 s 4526 39200 4582 40000 0 FreeSans 224 90 0 0 s_wb_adr[1]
port 83 nsew signal tristate
flabel metal2 s 15014 39200 15070 40000 0 FreeSans 224 90 0 0 s_wb_adr[20]
port 84 nsew signal tristate
flabel metal2 s 15566 39200 15622 40000 0 FreeSans 224 90 0 0 s_wb_adr[21]
port 85 nsew signal tristate
flabel metal2 s 16118 39200 16174 40000 0 FreeSans 224 90 0 0 s_wb_adr[22]
port 86 nsew signal tristate
flabel metal2 s 16670 39200 16726 40000 0 FreeSans 224 90 0 0 s_wb_adr[23]
port 87 nsew signal tristate
flabel metal2 s 5078 39200 5134 40000 0 FreeSans 224 90 0 0 s_wb_adr[2]
port 88 nsew signal tristate
flabel metal2 s 5630 39200 5686 40000 0 FreeSans 224 90 0 0 s_wb_adr[3]
port 89 nsew signal tristate
flabel metal2 s 6182 39200 6238 40000 0 FreeSans 224 90 0 0 s_wb_adr[4]
port 90 nsew signal tristate
flabel metal2 s 6734 39200 6790 40000 0 FreeSans 224 90 0 0 s_wb_adr[5]
port 91 nsew signal tristate
flabel metal2 s 7286 39200 7342 40000 0 FreeSans 224 90 0 0 s_wb_adr[6]
port 92 nsew signal tristate
flabel metal2 s 7838 39200 7894 40000 0 FreeSans 224 90 0 0 s_wb_adr[7]
port 93 nsew signal tristate
flabel metal2 s 8390 39200 8446 40000 0 FreeSans 224 90 0 0 s_wb_adr[8]
port 94 nsew signal tristate
flabel metal2 s 8942 39200 8998 40000 0 FreeSans 224 90 0 0 s_wb_adr[9]
port 95 nsew signal tristate
flabel metal2 s 17222 39200 17278 40000 0 FreeSans 224 90 0 0 s_wb_cyc
port 96 nsew signal tristate
flabel metal2 s 17774 39200 17830 40000 0 FreeSans 224 90 0 0 s_wb_err
port 97 nsew signal input
flabel metal2 s 18326 39200 18382 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[0]
port 98 nsew signal input
flabel metal2 s 23846 39200 23902 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[10]
port 99 nsew signal input
flabel metal2 s 24398 39200 24454 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[11]
port 100 nsew signal input
flabel metal2 s 24950 39200 25006 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[12]
port 101 nsew signal input
flabel metal2 s 25502 39200 25558 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[13]
port 102 nsew signal input
flabel metal2 s 26054 39200 26110 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[14]
port 103 nsew signal input
flabel metal2 s 26606 39200 26662 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[15]
port 104 nsew signal input
flabel metal2 s 18878 39200 18934 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[1]
port 105 nsew signal input
flabel metal2 s 19430 39200 19486 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[2]
port 106 nsew signal input
flabel metal2 s 19982 39200 20038 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[3]
port 107 nsew signal input
flabel metal2 s 20534 39200 20590 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[4]
port 108 nsew signal input
flabel metal2 s 21086 39200 21142 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[5]
port 109 nsew signal input
flabel metal2 s 21638 39200 21694 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[6]
port 110 nsew signal input
flabel metal2 s 22190 39200 22246 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[7]
port 111 nsew signal input
flabel metal2 s 22742 39200 22798 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[8]
port 112 nsew signal input
flabel metal2 s 23294 39200 23350 40000 0 FreeSans 224 90 0 0 s_wb_i_dat[9]
port 113 nsew signal input
flabel metal2 s 27158 39200 27214 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[0]
port 114 nsew signal tristate
flabel metal2 s 32678 39200 32734 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[10]
port 115 nsew signal tristate
flabel metal2 s 33230 39200 33286 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[11]
port 116 nsew signal tristate
flabel metal2 s 33782 39200 33838 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[12]
port 117 nsew signal tristate
flabel metal2 s 34334 39200 34390 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[13]
port 118 nsew signal tristate
flabel metal2 s 34886 39200 34942 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[14]
port 119 nsew signal tristate
flabel metal2 s 35438 39200 35494 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[15]
port 120 nsew signal tristate
flabel metal2 s 27710 39200 27766 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[1]
port 121 nsew signal tristate
flabel metal2 s 28262 39200 28318 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[2]
port 122 nsew signal tristate
flabel metal2 s 28814 39200 28870 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[3]
port 123 nsew signal tristate
flabel metal2 s 29366 39200 29422 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[4]
port 124 nsew signal tristate
flabel metal2 s 29918 39200 29974 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[5]
port 125 nsew signal tristate
flabel metal2 s 30470 39200 30526 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[6]
port 126 nsew signal tristate
flabel metal2 s 31022 39200 31078 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[7]
port 127 nsew signal tristate
flabel metal2 s 31574 39200 31630 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[8]
port 128 nsew signal tristate
flabel metal2 s 32126 39200 32182 40000 0 FreeSans 224 90 0 0 s_wb_o_dat[9]
port 129 nsew signal tristate
flabel metal2 s 35990 39200 36046 40000 0 FreeSans 224 90 0 0 s_wb_sel[0]
port 130 nsew signal tristate
flabel metal2 s 36542 39200 36598 40000 0 FreeSans 224 90 0 0 s_wb_sel[1]
port 131 nsew signal tristate
flabel metal2 s 37094 39200 37150 40000 0 FreeSans 224 90 0 0 s_wb_stb
port 132 nsew signal tristate
flabel metal2 s 37646 39200 37702 40000 0 FreeSans 224 90 0 0 s_wb_we
port 133 nsew signal tristate
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 134 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 134 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 135 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
